-- Generated from Simulink block PSB3_0/0001_
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_0001 is
  port (
    rst : in std_logic_vector( 1-1 downto 0 );
    en : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    out_x0 : out std_logic_vector( 1-1 downto 0 )
  );
end psb3_0_0001;
architecture structural of psb3_0_0001 is 
  signal gin_tl_reset_net : std_logic_vector( 1-1 downto 0 );
  signal constant17_op_net : std_logic_vector( 2-1 downto 0 );
  signal register_q_net : std_logic_vector( 1-1 downto 0 );
  signal gin_tl_start_net : std_logic_vector( 1-1 downto 0 );
  signal counter_op_net : std_logic_vector( 2-1 downto 0 );
  signal const_op_net : std_logic_vector( 1-1 downto 0 );
  signal relational_op_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal ce_net : std_logic;
begin
  out_x0 <= register_q_net;
  gin_tl_reset_net <= rst;
  gin_tl_start_net <= en;
  clk_net <= clk_1;
  ce_net <= ce_1;
  constant17 : entity xil_defaultlib.sysgen_constant_e0cdecfe1b 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant17_op_net
  );
  counter : entity xil_defaultlib.psb3_0_xlcounter_free 
  generic map (
    core_name0 => "psb3_0_c_counter_binary_v12_0_i1",
    op_arith => xlUnsigned,
    op_width => 2
  )
  port map (
    clr => '0',
    rst => gin_tl_reset_net,
    en => gin_tl_start_net,
    clk => clk_net,
    ce => ce_net,
    op => counter_op_net
  );
  register_x0 : entity xil_defaultlib.psb3_0_xlregister 
  generic map (
    d_width => 1,
    init_value => b"0"
  )
  port map (
    d => const_op_net,
    rst => gin_tl_reset_net,
    en => relational_op_net,
    clk => clk_net,
    ce => ce_net,
    q => register_q_net
  );
  relational : entity xil_defaultlib.sysgen_relational_499eab296f 
  port map (
    clr => '0',
    a => counter_op_net,
    b => constant17_op_net,
    clk => clk_net,
    ce => ce_net,
    op => relational_op_net
  );
  const : entity xil_defaultlib.sysgen_constant_71e89d757c 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => const_op_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Baseband_even_1/delayCounter2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_delaycounter2 is
  port (
    edge1 : in std_logic_vector( 1-1 downto 0 );
    edge2 : in std_logic;
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    delay : out std_logic_vector( 12-1 downto 0 )
  );
end psb3_0_delaycounter2;
architecture structural of psb3_0_delaycounter2 is 
  signal ce_net : std_logic;
  signal register1_q_net : std_logic_vector( 1-1 downto 0 );
  signal register2_q_net : std_logic_vector( 1-1 downto 0 );
  signal counter1_op_net : std_logic_vector( 12-1 downto 0 );
  signal delay14_q_net : std_logic_vector( 1-1 downto 0 );
  signal cordic_6_0_even_1_m_axis_dout_tvalid_net : std_logic;
  signal clk_net : std_logic;
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
  signal const1_op_net : std_logic_vector( 1-1 downto 0 );
begin
  delay <= counter1_op_net;
  delay14_q_net <= edge1;
  cordic_6_0_even_1_m_axis_dout_tvalid_net <= edge2;
  clk_net <= clk_1;
  ce_net <= ce_1;
  counter1 : entity xil_defaultlib.psb3_0_xlcounter_free 
  generic map (
    core_name0 => "psb3_0_c_counter_binary_v12_0_i2",
    op_arith => xlUnsigned,
    op_width => 12
  )
  port map (
    rst => "0",
    clr => '0',
    en => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    op => counter1_op_net
  );
  logical : entity xil_defaultlib.sysgen_logical_e072b658e1 
  port map (
    clr => '0',
    d0 => register1_q_net,
    d1 => register2_q_net,
    clk => clk_net,
    ce => ce_net,
    y => logical_y_net
  );
  register1 : entity xil_defaultlib.psb3_0_xlregister 
  generic map (
    d_width => 1,
    init_value => b"0"
  )
  port map (
    rst => "0",
    d => const1_op_net,
    en => delay14_q_net,
    clk => clk_net,
    ce => ce_net,
    q => register1_q_net
  );
  register2 : entity xil_defaultlib.psb3_0_xlregister 
  generic map (
    d_width => 1,
    init_value => b"0"
  )
  port map (
    rst => "0",
    d => const1_op_net,
    en(0) => cordic_6_0_even_1_m_axis_dout_tvalid_net,
    clk => clk_net,
    ce => ce_net,
    q => register2_q_net
  );
  const1 : entity xil_defaultlib.sysgen_constant_71e89d757c 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => const1_op_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Baseband_even_1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_baseband_even_1 is
  port (
    in_tvalid : in std_logic_vector( 1-1 downto 0 );
    addr_r : in std_logic_vector( 8-1 downto 0 );
    addr_w : in std_logic_vector( 8-1 downto 0 );
    init_im_even : in std_logic_vector( 18-1 downto 0 );
    init_re_even : in std_logic_vector( 18-1 downto 0 );
    dphi_even : in std_logic_vector( 16-1 downto 0 );
    we : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    delay_count : out std_logic_vector( 12-1 downto 0 );
    out_im : out std_logic_vector( 16-1 downto 0 );
    out_re : out std_logic_vector( 16-1 downto 0 );
    out_tvalid : out std_logic
  );
end psb3_0_baseband_even_1;
architecture structural of psb3_0_baseband_even_1 is 
  signal dpram_dphi_even_1_douta_net : std_logic_vector( 16-1 downto 0 );
  signal delay37_q_net : std_logic_vector( 16-1 downto 0 );
  signal delay35_q_net : std_logic_vector( 18-1 downto 0 );
  signal cordic_6_0_even_1_m_axis_dout_tdata_real_net : std_logic_vector( 16-1 downto 0 );
  signal ram_dphi_addr_op_net : std_logic_vector( 8-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal ce_net : std_logic;
  signal delay14_q_net : std_logic_vector( 1-1 downto 0 );
  signal counter1_op_net : std_logic_vector( 12-1 downto 0 );
  signal addsub_s_net : std_logic_vector( 16-1 downto 0 );
  signal fifo4_dout_net : std_logic_vector( 16-1 downto 0 );
  signal cordic_6_0_even_1_m_axis_dout_tvalid_net : std_logic;
  signal cordic_6_0_even_1_m_axis_dout_tdata_imag_net : std_logic_vector( 16-1 downto 0 );
  signal delay38_q_net : std_logic_vector( 8-1 downto 0 );
  signal delay44_q_net : std_logic_vector( 18-1 downto 0 );
  signal constant7_op_net : std_logic_vector( 18-1 downto 0 );
  signal constant2_op_net : std_logic_vector( 1-1 downto 0 );
  signal constant_op_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal constant8_op_net : std_logic_vector( 16-1 downto 0 );
  signal dpram_init_im_even_1_douta_net : std_logic_vector( 18-1 downto 0 );
  signal dpram_init_re_even_1_douta_net : std_logic_vector( 18-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 1-1 downto 0 );
  signal constant6_op_net : std_logic_vector( 1-1 downto 0 );
  signal convert2_dout_net : std_logic_vector( 18-1 downto 0 );
  signal constant3_op_net : std_logic_vector( 18-1 downto 0 );
  signal dpram_init_re_even_1_doutb_net : std_logic_vector( 18-1 downto 0 );
  signal dpram_dphi_even_1_doutb_net : std_logic_vector( 16-1 downto 0 );
  signal delay16_q_net : std_logic_vector( 1-1 downto 0 );
  signal fifo4_empty_net : std_logic;
  signal fifo4_full_net : std_logic;
  signal dpram_init_im_even_1_doutb_net : std_logic_vector( 18-1 downto 0 );
begin
  delay_count <= counter1_op_net;
  out_im <= cordic_6_0_even_1_m_axis_dout_tdata_imag_net;
  out_re <= cordic_6_0_even_1_m_axis_dout_tdata_real_net;
  out_tvalid <= cordic_6_0_even_1_m_axis_dout_tvalid_net;
  delay14_q_net <= in_tvalid;
  ram_dphi_addr_op_net <= addr_r;
  delay38_q_net <= addr_w;
  delay44_q_net <= init_im_even;
  delay35_q_net <= init_re_even;
  delay37_q_net <= dphi_even;
  delay1_q_net <= we;
  clk_net <= clk_1;
  ce_net <= ce_1;
  delaycounter2_x0 : entity xil_defaultlib.psb3_0_delaycounter2 
  port map (
    edge1 => delay14_q_net,
    edge2 => cordic_6_0_even_1_m_axis_dout_tvalid_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    delay => counter1_op_net
  );
  addsub : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 16,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 17,
    core_name0 => "psb3_0_c_addsub_v12_0_i0",
    extra_registers => 1,
    full_s_arith => 1,
    full_s_width => 17,
    latency => 2,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => dpram_dphi_even_1_douta_net,
    b => fifo4_dout_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  cordic_6_0_even_1 : entity xil_defaultlib.xlcordic_5a76bbdd6458ef1eb96e9ff32fab9279 
  port map (
    s_axis_cartesian_tvalid => delay14_q_net(0),
    s_axis_cartesian_tdata_imag => dpram_init_im_even_1_douta_net,
    s_axis_cartesian_tdata_real => dpram_init_re_even_1_douta_net,
    s_axis_phase_tvalid => delay14_q_net(0),
    s_axis_phase_tdata_phase => convert2_dout_net,
    clk => clk_net,
    ce => ce_net,
    m_axis_dout_tvalid => cordic_6_0_even_1_m_axis_dout_tvalid_net,
    m_axis_dout_tdata_imag => cordic_6_0_even_1_m_axis_dout_tdata_imag_net,
    m_axis_dout_tdata_real => cordic_6_0_even_1_m_axis_dout_tdata_real_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_de9059c03f 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_de9059c03f 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  constant2 : entity xil_defaultlib.sysgen_constant_de9059c03f 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant2_op_net
  );
  constant3 : entity xil_defaultlib.sysgen_constant_ac4aa5284f 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant3_op_net
  );
  constant6 : entity xil_defaultlib.sysgen_constant_71e89d757c 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant6_op_net
  );
  constant7 : entity xil_defaultlib.sysgen_constant_ac4aa5284f 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant7_op_net
  );
  constant8 : entity xil_defaultlib.sysgen_constant_eb74b92b90 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant8_op_net
  );
  convert2 : entity xil_defaultlib.psb3_0_xlconvert 
  generic map (
    bool_conversion => 0,
    din_arith => 2,
    din_bin_pt => 15,
    din_width => 16,
    dout_arith => 2,
    dout_bin_pt => 15,
    dout_width => 18,
    latency => 0,
    overflow => xlWrap,
    quantization => xlTruncate
  )
  port map (
    clr => '0',
    en => "1",
    din => reinterpret2_output_port_net,
    clk => clk_net,
    ce => ce_net,
    dout => convert2_dout_net
  );
  dpram_dphi_even_1 : entity xil_defaultlib.psb3_0_xltdpram 
  generic map (
    addr_width_b => 8,
    clocking_mode => "common_clock",
    data_width_b => 16,
    latency => 1,
    mem_init_file => "xpm_62c937_vivado.mem",
    mem_size => 4096,
    mem_type => "block",
    read_reset_a => "0",
    read_reset_b => "0",
    width => 16,
    width_addr => 8,
    write_mode_a => "read_first",
    write_mode_b => "read_first"
  )
  port map (
    ena => "1",
    enb => "1",
    rsta => "0",
    rstb => "0",
    addra => ram_dphi_addr_op_net,
    dina => constant8_op_net,
    wea => constant2_op_net,
    addrb => delay38_q_net,
    dinb => delay37_q_net,
    web => delay1_q_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dpram_dphi_even_1_douta_net,
    doutb => dpram_dphi_even_1_doutb_net
  );
  dpram_init_im_even_1 : entity xil_defaultlib.psb3_0_xltdpram 
  generic map (
    addr_width_b => 8,
    clocking_mode => "common_clock",
    data_width_b => 18,
    latency => 1,
    mem_init_file => "xpm_c13bdd_vivado.mem",
    mem_size => 4608,
    mem_type => "block",
    read_reset_a => "0",
    read_reset_b => "0",
    width => 18,
    width_addr => 8,
    write_mode_a => "read_first",
    write_mode_b => "read_first"
  )
  port map (
    ena => "1",
    enb => "1",
    rsta => "0",
    rstb => "0",
    addra => ram_dphi_addr_op_net,
    dina => constant3_op_net,
    wea => constant_op_net,
    addrb => delay38_q_net,
    dinb => delay44_q_net,
    web => delay1_q_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dpram_init_im_even_1_douta_net,
    doutb => dpram_init_im_even_1_doutb_net
  );
  dpram_init_re_even_1 : entity xil_defaultlib.psb3_0_xltdpram 
  generic map (
    addr_width_b => 8,
    clocking_mode => "common_clock",
    data_width_b => 18,
    latency => 1,
    mem_init_file => "xpm_26a6e7_vivado.mem",
    mem_size => 4608,
    mem_type => "block",
    read_reset_a => "0",
    read_reset_b => "0",
    width => 18,
    width_addr => 8,
    write_mode_a => "read_first",
    write_mode_b => "read_first"
  )
  port map (
    ena => "1",
    enb => "1",
    rsta => "0",
    rstb => "0",
    addra => ram_dphi_addr_op_net,
    dina => constant7_op_net,
    wea => constant1_op_net,
    addrb => delay38_q_net,
    dinb => delay35_q_net,
    web => delay1_q_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dpram_init_re_even_1_douta_net,
    doutb => dpram_init_re_even_1_doutb_net
  );
  delay16 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 253,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => constant6_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay16_q_net
  );
  fifo4 : entity xil_defaultlib.psb3_0_xlfifogen_u 
  generic map (
    core_name0 => "psb3_0_fifo_generator_i1",
    data_count_width => 10,
    data_width => 16,
    extra_registers => 1,
    has_ae => 0,
    has_af => 0,
    has_rst => false,
    ignore_din_for_gcd => false,
    percent_full_width => 1
  )
  port map (
    en => '1',
    rst => '0',
    din => addsub_s_net,
    we => constant6_op_net(0),
    re => delay16_q_net(0),
    clk => clk_net,
    ce => ce_net,
    we_ce => ce_net,
    re_ce => ce_net,
    dout => fifo4_dout_net,
    empty => fifo4_empty_net,
    full => fifo4_full_net
  );
  reinterpret2 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => fifo4_dout_net,
    output_port => reinterpret2_output_port_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Baseband_even_2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_baseband_even_2 is
  port (
    in_tvalid : in std_logic_vector( 1-1 downto 0 );
    addr_r : in std_logic_vector( 8-1 downto 0 );
    addr_w : in std_logic_vector( 8-1 downto 0 );
    init_im_even_2 : in std_logic_vector( 18-1 downto 0 );
    init_re_even_2 : in std_logic_vector( 18-1 downto 0 );
    dphi_even_2 : in std_logic_vector( 16-1 downto 0 );
    we : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    out_im : out std_logic_vector( 16-1 downto 0 );
    out_re : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_baseband_even_2;
architecture structural of psb3_0_baseband_even_2 is 
  signal delay37_q_net : std_logic_vector( 16-1 downto 0 );
  signal dpram_dphi_even_2_douta_net : std_logic_vector( 16-1 downto 0 );
  signal cordic_6_0_even_2_m_axis_dout_tdata_imag_net : std_logic_vector( 16-1 downto 0 );
  signal convert2_dout_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal cordic_6_0_even_2_m_axis_dout_tvalid_net : std_logic;
  signal cordic_6_0_even_2_m_axis_dout_tdata_real_net : std_logic_vector( 16-1 downto 0 );
  signal dpram_init_im_even_2_douta_net : std_logic_vector( 18-1 downto 0 );
  signal delay35_q_net : std_logic_vector( 18-1 downto 0 );
  signal ram_dphi_addr_op_net : std_logic_vector( 8-1 downto 0 );
  signal delay14_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay44_q_net : std_logic_vector( 18-1 downto 0 );
  signal fifo4_dout_net : std_logic_vector( 16-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 1-1 downto 0 );
  signal addsub_s_net : std_logic_vector( 16-1 downto 0 );
  signal delay38_q_net : std_logic_vector( 8-1 downto 0 );
  signal ce_net : std_logic;
  signal dpram_init_re_even_2_douta_net : std_logic_vector( 18-1 downto 0 );
  signal constant_op_net : std_logic_vector( 1-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 1-1 downto 0 );
  signal constant2_op_net : std_logic_vector( 1-1 downto 0 );
  signal constant6_op_net : std_logic_vector( 1-1 downto 0 );
  signal dpram_dphi_even_2_doutb_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal constant7_op_net : std_logic_vector( 18-1 downto 0 );
  signal constant8_op_net : std_logic_vector( 16-1 downto 0 );
  signal constant3_op_net : std_logic_vector( 18-1 downto 0 );
  signal delay16_q_net : std_logic_vector( 1-1 downto 0 );
  signal dpram_init_re_even_2_doutb_net : std_logic_vector( 18-1 downto 0 );
  signal dpram_init_im_even_2_doutb_net : std_logic_vector( 18-1 downto 0 );
  signal fifo4_empty_net : std_logic;
  signal fifo4_full_net : std_logic;
begin
  out_im <= cordic_6_0_even_2_m_axis_dout_tdata_imag_net;
  out_re <= cordic_6_0_even_2_m_axis_dout_tdata_real_net;
  delay14_q_net <= in_tvalid;
  ram_dphi_addr_op_net <= addr_r;
  delay38_q_net <= addr_w;
  delay44_q_net <= init_im_even_2;
  delay35_q_net <= init_re_even_2;
  delay37_q_net <= dphi_even_2;
  delay8_q_net <= we;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 16,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 17,
    core_name0 => "psb3_0_c_addsub_v12_0_i0",
    extra_registers => 1,
    full_s_arith => 1,
    full_s_width => 17,
    latency => 2,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => dpram_dphi_even_2_douta_net,
    b => fifo4_dout_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  cordic_6_0_even_2 : entity xil_defaultlib.xlcordic_5a76bbdd6458ef1eb96e9ff32fab9279 
  port map (
    s_axis_cartesian_tvalid => delay14_q_net(0),
    s_axis_cartesian_tdata_imag => dpram_init_im_even_2_douta_net,
    s_axis_cartesian_tdata_real => dpram_init_re_even_2_douta_net,
    s_axis_phase_tvalid => delay14_q_net(0),
    s_axis_phase_tdata_phase => convert2_dout_net,
    clk => clk_net,
    ce => ce_net,
    m_axis_dout_tvalid => cordic_6_0_even_2_m_axis_dout_tvalid_net,
    m_axis_dout_tdata_imag => cordic_6_0_even_2_m_axis_dout_tdata_imag_net,
    m_axis_dout_tdata_real => cordic_6_0_even_2_m_axis_dout_tdata_real_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_de9059c03f 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_de9059c03f 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  constant2 : entity xil_defaultlib.sysgen_constant_de9059c03f 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant2_op_net
  );
  constant3 : entity xil_defaultlib.sysgen_constant_ac4aa5284f 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant3_op_net
  );
  constant6 : entity xil_defaultlib.sysgen_constant_71e89d757c 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant6_op_net
  );
  constant7 : entity xil_defaultlib.sysgen_constant_ac4aa5284f 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant7_op_net
  );
  constant8 : entity xil_defaultlib.sysgen_constant_eb74b92b90 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant8_op_net
  );
  convert2 : entity xil_defaultlib.psb3_0_xlconvert 
  generic map (
    bool_conversion => 0,
    din_arith => 2,
    din_bin_pt => 15,
    din_width => 16,
    dout_arith => 2,
    dout_bin_pt => 15,
    dout_width => 18,
    latency => 0,
    overflow => xlWrap,
    quantization => xlTruncate
  )
  port map (
    clr => '0',
    en => "1",
    din => reinterpret2_output_port_net,
    clk => clk_net,
    ce => ce_net,
    dout => convert2_dout_net
  );
  dpram_dphi_even_2 : entity xil_defaultlib.psb3_0_xltdpram 
  generic map (
    addr_width_b => 8,
    clocking_mode => "common_clock",
    data_width_b => 16,
    latency => 1,
    mem_init_file => "xpm_908ac5_vivado.mem",
    mem_size => 4096,
    mem_type => "block",
    read_reset_a => "0",
    read_reset_b => "0",
    width => 16,
    width_addr => 8,
    write_mode_a => "read_first",
    write_mode_b => "read_first"
  )
  port map (
    ena => "1",
    enb => "1",
    rsta => "0",
    rstb => "0",
    addra => ram_dphi_addr_op_net,
    dina => constant8_op_net,
    wea => constant2_op_net,
    addrb => delay38_q_net,
    dinb => delay37_q_net,
    web => delay8_q_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dpram_dphi_even_2_douta_net,
    doutb => dpram_dphi_even_2_doutb_net
  );
  dpram_init_im_even_2 : entity xil_defaultlib.psb3_0_xltdpram 
  generic map (
    addr_width_b => 8,
    clocking_mode => "common_clock",
    data_width_b => 18,
    latency => 1,
    mem_init_file => "xpm_3d0358_vivado.mem",
    mem_size => 4608,
    mem_type => "block",
    read_reset_a => "0",
    read_reset_b => "0",
    width => 18,
    width_addr => 8,
    write_mode_a => "read_first",
    write_mode_b => "read_first"
  )
  port map (
    ena => "1",
    enb => "1",
    rsta => "0",
    rstb => "0",
    addra => ram_dphi_addr_op_net,
    dina => constant3_op_net,
    wea => constant_op_net,
    addrb => delay38_q_net,
    dinb => delay44_q_net,
    web => delay8_q_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dpram_init_im_even_2_douta_net,
    doutb => dpram_init_im_even_2_doutb_net
  );
  dpram_init_re_even_2 : entity xil_defaultlib.psb3_0_xltdpram 
  generic map (
    addr_width_b => 8,
    clocking_mode => "common_clock",
    data_width_b => 18,
    latency => 1,
    mem_init_file => "xpm_20e520_vivado.mem",
    mem_size => 4608,
    mem_type => "block",
    read_reset_a => "0",
    read_reset_b => "0",
    width => 18,
    width_addr => 8,
    write_mode_a => "read_first",
    write_mode_b => "read_first"
  )
  port map (
    ena => "1",
    enb => "1",
    rsta => "0",
    rstb => "0",
    addra => ram_dphi_addr_op_net,
    dina => constant7_op_net,
    wea => constant1_op_net,
    addrb => delay38_q_net,
    dinb => delay35_q_net,
    web => delay8_q_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dpram_init_re_even_2_douta_net,
    doutb => dpram_init_re_even_2_doutb_net
  );
  delay16 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 253,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => constant6_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay16_q_net
  );
  fifo4 : entity xil_defaultlib.psb3_0_xlfifogen_u 
  generic map (
    core_name0 => "psb3_0_fifo_generator_i1",
    data_count_width => 10,
    data_width => 16,
    extra_registers => 1,
    has_ae => 0,
    has_af => 0,
    has_rst => false,
    ignore_din_for_gcd => false,
    percent_full_width => 1
  )
  port map (
    en => '1',
    rst => '0',
    din => addsub_s_net,
    we => constant6_op_net(0),
    re => delay16_q_net(0),
    clk => clk_net,
    ce => ce_net,
    we_ce => ce_net,
    re_ce => ce_net,
    dout => fifo4_dout_net,
    empty => fifo4_empty_net,
    full => fifo4_full_net
  );
  reinterpret2 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => fifo4_dout_net,
    output_port => reinterpret2_output_port_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Baseband_even_3
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_baseband_even_3 is
  port (
    in_tvalid : in std_logic_vector( 1-1 downto 0 );
    addr_r : in std_logic_vector( 8-1 downto 0 );
    addr_w : in std_logic_vector( 8-1 downto 0 );
    init_im_even : in std_logic_vector( 18-1 downto 0 );
    init_re_even : in std_logic_vector( 18-1 downto 0 );
    dphi_even : in std_logic_vector( 16-1 downto 0 );
    we : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    out_im : out std_logic_vector( 16-1 downto 0 );
    out_re : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_baseband_even_3;
architecture structural of psb3_0_baseband_even_3 is 
  signal constant8_op_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal dpram_dphi_even_3_doutb_net : std_logic_vector( 16-1 downto 0 );
  signal dpram_init_re_even_3_doutb_net : std_logic_vector( 18-1 downto 0 );
  signal dpram_init_im_even_3_doutb_net : std_logic_vector( 18-1 downto 0 );
  signal delay16_q_net : std_logic_vector( 1-1 downto 0 );
  signal fifo4_empty_net : std_logic;
  signal fifo4_full_net : std_logic;
  signal constant_op_net : std_logic_vector( 1-1 downto 0 );
  signal constant2_op_net : std_logic_vector( 1-1 downto 0 );
  signal dpram_init_im_even_3_douta_net : std_logic_vector( 18-1 downto 0 );
  signal fifo4_dout_net : std_logic_vector( 16-1 downto 0 );
  signal constant3_op_net : std_logic_vector( 18-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 1-1 downto 0 );
  signal cordic_6_0_even_1_m_axis_dout_tvalid_net : std_logic;
  signal dpram_init_re_even_3_douta_net : std_logic_vector( 18-1 downto 0 );
  signal dpram_dphi_even_3_douta_net : std_logic_vector( 16-1 downto 0 );
  signal constant6_op_net : std_logic_vector( 1-1 downto 0 );
  signal constant7_op_net : std_logic_vector( 18-1 downto 0 );
  signal addsub_s_net : std_logic_vector( 16-1 downto 0 );
  signal convert2_dout_net : std_logic_vector( 18-1 downto 0 );
  signal cordic_6_0_even_1_m_axis_dout_tdata_imag_net : std_logic_vector( 16-1 downto 0 );
  signal delay44_q_net : std_logic_vector( 18-1 downto 0 );
  signal ram_dphi_addr_op_net : std_logic_vector( 8-1 downto 0 );
  signal cordic_6_0_even_1_m_axis_dout_tdata_real_net : std_logic_vector( 16-1 downto 0 );
  signal delay14_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay38_q_net : std_logic_vector( 8-1 downto 0 );
  signal delay35_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay37_q_net : std_logic_vector( 16-1 downto 0 );
  signal delay31_q_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal ce_net : std_logic;
begin
  out_im <= cordic_6_0_even_1_m_axis_dout_tdata_imag_net;
  out_re <= cordic_6_0_even_1_m_axis_dout_tdata_real_net;
  delay14_q_net <= in_tvalid;
  ram_dphi_addr_op_net <= addr_r;
  delay38_q_net <= addr_w;
  delay44_q_net <= init_im_even;
  delay35_q_net <= init_re_even;
  delay37_q_net <= dphi_even;
  delay31_q_net <= we;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 16,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 17,
    core_name0 => "psb3_0_c_addsub_v12_0_i0",
    extra_registers => 1,
    full_s_arith => 1,
    full_s_width => 17,
    latency => 2,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => dpram_dphi_even_3_douta_net,
    b => fifo4_dout_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  cordic_6_0_even_1 : entity xil_defaultlib.xlcordic_5a76bbdd6458ef1eb96e9ff32fab9279 
  port map (
    s_axis_cartesian_tvalid => delay14_q_net(0),
    s_axis_cartesian_tdata_imag => dpram_init_im_even_3_douta_net,
    s_axis_cartesian_tdata_real => dpram_init_re_even_3_douta_net,
    s_axis_phase_tvalid => delay14_q_net(0),
    s_axis_phase_tdata_phase => convert2_dout_net,
    clk => clk_net,
    ce => ce_net,
    m_axis_dout_tvalid => cordic_6_0_even_1_m_axis_dout_tvalid_net,
    m_axis_dout_tdata_imag => cordic_6_0_even_1_m_axis_dout_tdata_imag_net,
    m_axis_dout_tdata_real => cordic_6_0_even_1_m_axis_dout_tdata_real_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_de9059c03f 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_de9059c03f 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  constant2 : entity xil_defaultlib.sysgen_constant_de9059c03f 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant2_op_net
  );
  constant3 : entity xil_defaultlib.sysgen_constant_ac4aa5284f 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant3_op_net
  );
  constant6 : entity xil_defaultlib.sysgen_constant_71e89d757c 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant6_op_net
  );
  constant7 : entity xil_defaultlib.sysgen_constant_ac4aa5284f 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant7_op_net
  );
  constant8 : entity xil_defaultlib.sysgen_constant_eb74b92b90 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant8_op_net
  );
  convert2 : entity xil_defaultlib.psb3_0_xlconvert 
  generic map (
    bool_conversion => 0,
    din_arith => 2,
    din_bin_pt => 15,
    din_width => 16,
    dout_arith => 2,
    dout_bin_pt => 15,
    dout_width => 18,
    latency => 0,
    overflow => xlWrap,
    quantization => xlTruncate
  )
  port map (
    clr => '0',
    en => "1",
    din => reinterpret2_output_port_net,
    clk => clk_net,
    ce => ce_net,
    dout => convert2_dout_net
  );
  dpram_dphi_even_3 : entity xil_defaultlib.psb3_0_xltdpram 
  generic map (
    addr_width_b => 8,
    clocking_mode => "common_clock",
    data_width_b => 16,
    latency => 1,
    mem_init_file => "xpm_9a918a_vivado.mem",
    mem_size => 4096,
    mem_type => "block",
    read_reset_a => "0",
    read_reset_b => "0",
    width => 16,
    width_addr => 8,
    write_mode_a => "read_first",
    write_mode_b => "read_first"
  )
  port map (
    ena => "1",
    enb => "1",
    rsta => "0",
    rstb => "0",
    addra => ram_dphi_addr_op_net,
    dina => constant8_op_net,
    wea => constant2_op_net,
    addrb => delay38_q_net,
    dinb => delay37_q_net,
    web => delay31_q_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dpram_dphi_even_3_douta_net,
    doutb => dpram_dphi_even_3_doutb_net
  );
  dpram_init_im_even_3 : entity xil_defaultlib.psb3_0_xltdpram 
  generic map (
    addr_width_b => 8,
    clocking_mode => "common_clock",
    data_width_b => 18,
    latency => 1,
    mem_init_file => "xpm_1f4a12_vivado.mem",
    mem_size => 4608,
    mem_type => "block",
    read_reset_a => "0",
    read_reset_b => "0",
    width => 18,
    width_addr => 8,
    write_mode_a => "read_first",
    write_mode_b => "read_first"
  )
  port map (
    ena => "1",
    enb => "1",
    rsta => "0",
    rstb => "0",
    addra => ram_dphi_addr_op_net,
    dina => constant3_op_net,
    wea => constant_op_net,
    addrb => delay38_q_net,
    dinb => delay44_q_net,
    web => delay31_q_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dpram_init_im_even_3_douta_net,
    doutb => dpram_init_im_even_3_doutb_net
  );
  dpram_init_re_even_3 : entity xil_defaultlib.psb3_0_xltdpram 
  generic map (
    addr_width_b => 8,
    clocking_mode => "common_clock",
    data_width_b => 18,
    latency => 1,
    mem_init_file => "xpm_6d9a13_vivado.mem",
    mem_size => 4608,
    mem_type => "block",
    read_reset_a => "0",
    read_reset_b => "0",
    width => 18,
    width_addr => 8,
    write_mode_a => "read_first",
    write_mode_b => "read_first"
  )
  port map (
    ena => "1",
    enb => "1",
    rsta => "0",
    rstb => "0",
    addra => ram_dphi_addr_op_net,
    dina => constant7_op_net,
    wea => constant1_op_net,
    addrb => delay38_q_net,
    dinb => delay35_q_net,
    web => delay31_q_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dpram_init_re_even_3_douta_net,
    doutb => dpram_init_re_even_3_doutb_net
  );
  delay16 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 253,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => constant6_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay16_q_net
  );
  fifo4 : entity xil_defaultlib.psb3_0_xlfifogen_u 
  generic map (
    core_name0 => "psb3_0_fifo_generator_i1",
    data_count_width => 10,
    data_width => 16,
    extra_registers => 1,
    has_ae => 0,
    has_af => 0,
    has_rst => false,
    ignore_din_for_gcd => false,
    percent_full_width => 1
  )
  port map (
    en => '1',
    rst => '0',
    din => addsub_s_net,
    we => constant6_op_net(0),
    re => delay16_q_net(0),
    clk => clk_net,
    ce => ce_net,
    we_ce => ce_net,
    re_ce => ce_net,
    dout => fifo4_dout_net,
    empty => fifo4_empty_net,
    full => fifo4_full_net
  );
  reinterpret2 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => fifo4_dout_net,
    output_port => reinterpret2_output_port_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Baseband_even_4
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_baseband_even_4 is
  port (
    in_tvalid : in std_logic_vector( 1-1 downto 0 );
    addr_r : in std_logic_vector( 8-1 downto 0 );
    addr_w : in std_logic_vector( 8-1 downto 0 );
    init_im_even_2 : in std_logic_vector( 18-1 downto 0 );
    init_re_even_2 : in std_logic_vector( 18-1 downto 0 );
    dphi_even_2 : in std_logic_vector( 16-1 downto 0 );
    we : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    out_im : out std_logic_vector( 16-1 downto 0 );
    out_re : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_baseband_even_4;
architecture structural of psb3_0_baseband_even_4 is 
  signal cordic_6_0_even_2_m_axis_dout_tdata_real_net : std_logic_vector( 16-1 downto 0 );
  signal delay14_q_net : std_logic_vector( 1-1 downto 0 );
  signal ram_dphi_addr_op_net : std_logic_vector( 8-1 downto 0 );
  signal delay38_q_net : std_logic_vector( 8-1 downto 0 );
  signal delay44_q_net : std_logic_vector( 18-1 downto 0 );
  signal cordic_6_0_even_2_m_axis_dout_tdata_imag_net : std_logic_vector( 16-1 downto 0 );
  signal delay49_q_net : std_logic_vector( 1-1 downto 0 );
  signal dpram_dphi_even_4_douta_net : std_logic_vector( 16-1 downto 0 );
  signal fifo4_dout_net : std_logic_vector( 16-1 downto 0 );
  signal clk_net : std_logic;
  signal cordic_6_0_even_2_m_axis_dout_tvalid_net : std_logic;
  signal dpram_init_im_even_4_douta_net : std_logic_vector( 18-1 downto 0 );
  signal dpram_init_re_even_4_douta_net : std_logic_vector( 18-1 downto 0 );
  signal delay35_q_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal addsub_s_net : std_logic_vector( 16-1 downto 0 );
  signal convert2_dout_net : std_logic_vector( 18-1 downto 0 );
  signal delay37_q_net : std_logic_vector( 16-1 downto 0 );
  signal constant2_op_net : std_logic_vector( 1-1 downto 0 );
  signal constant3_op_net : std_logic_vector( 18-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 1-1 downto 0 );
  signal constant7_op_net : std_logic_vector( 18-1 downto 0 );
  signal constant6_op_net : std_logic_vector( 1-1 downto 0 );
  signal constant_op_net : std_logic_vector( 1-1 downto 0 );
  signal constant8_op_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal dpram_dphi_even_4_doutb_net : std_logic_vector( 16-1 downto 0 );
  signal dpram_init_im_even_4_doutb_net : std_logic_vector( 18-1 downto 0 );
  signal dpram_init_re_even_4_doutb_net : std_logic_vector( 18-1 downto 0 );
  signal fifo4_empty_net : std_logic;
  signal delay16_q_net : std_logic_vector( 1-1 downto 0 );
  signal fifo4_full_net : std_logic;
begin
  out_im <= cordic_6_0_even_2_m_axis_dout_tdata_imag_net;
  out_re <= cordic_6_0_even_2_m_axis_dout_tdata_real_net;
  delay14_q_net <= in_tvalid;
  ram_dphi_addr_op_net <= addr_r;
  delay38_q_net <= addr_w;
  delay44_q_net <= init_im_even_2;
  delay35_q_net <= init_re_even_2;
  delay37_q_net <= dphi_even_2;
  delay49_q_net <= we;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 16,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 17,
    core_name0 => "psb3_0_c_addsub_v12_0_i0",
    extra_registers => 1,
    full_s_arith => 1,
    full_s_width => 17,
    latency => 2,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => dpram_dphi_even_4_douta_net,
    b => fifo4_dout_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  cordic_6_0_even_2 : entity xil_defaultlib.xlcordic_5a76bbdd6458ef1eb96e9ff32fab9279 
  port map (
    s_axis_cartesian_tvalid => delay14_q_net(0),
    s_axis_cartesian_tdata_imag => dpram_init_im_even_4_douta_net,
    s_axis_cartesian_tdata_real => dpram_init_re_even_4_douta_net,
    s_axis_phase_tvalid => delay14_q_net(0),
    s_axis_phase_tdata_phase => convert2_dout_net,
    clk => clk_net,
    ce => ce_net,
    m_axis_dout_tvalid => cordic_6_0_even_2_m_axis_dout_tvalid_net,
    m_axis_dout_tdata_imag => cordic_6_0_even_2_m_axis_dout_tdata_imag_net,
    m_axis_dout_tdata_real => cordic_6_0_even_2_m_axis_dout_tdata_real_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_de9059c03f 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_de9059c03f 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  constant2 : entity xil_defaultlib.sysgen_constant_de9059c03f 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant2_op_net
  );
  constant3 : entity xil_defaultlib.sysgen_constant_ac4aa5284f 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant3_op_net
  );
  constant6 : entity xil_defaultlib.sysgen_constant_71e89d757c 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant6_op_net
  );
  constant7 : entity xil_defaultlib.sysgen_constant_ac4aa5284f 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant7_op_net
  );
  constant8 : entity xil_defaultlib.sysgen_constant_eb74b92b90 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant8_op_net
  );
  convert2 : entity xil_defaultlib.psb3_0_xlconvert 
  generic map (
    bool_conversion => 0,
    din_arith => 2,
    din_bin_pt => 15,
    din_width => 16,
    dout_arith => 2,
    dout_bin_pt => 15,
    dout_width => 18,
    latency => 0,
    overflow => xlWrap,
    quantization => xlTruncate
  )
  port map (
    clr => '0',
    en => "1",
    din => reinterpret2_output_port_net,
    clk => clk_net,
    ce => ce_net,
    dout => convert2_dout_net
  );
  dpram_dphi_even_4 : entity xil_defaultlib.psb3_0_xltdpram 
  generic map (
    addr_width_b => 8,
    clocking_mode => "common_clock",
    data_width_b => 16,
    latency => 1,
    mem_init_file => "xpm_ec0e74_vivado.mem",
    mem_size => 4096,
    mem_type => "block",
    read_reset_a => "0",
    read_reset_b => "0",
    width => 16,
    width_addr => 8,
    write_mode_a => "read_first",
    write_mode_b => "read_first"
  )
  port map (
    ena => "1",
    enb => "1",
    rsta => "0",
    rstb => "0",
    addra => ram_dphi_addr_op_net,
    dina => constant8_op_net,
    wea => constant2_op_net,
    addrb => delay38_q_net,
    dinb => delay37_q_net,
    web => delay49_q_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dpram_dphi_even_4_douta_net,
    doutb => dpram_dphi_even_4_doutb_net
  );
  dpram_init_im_even_4 : entity xil_defaultlib.psb3_0_xltdpram 
  generic map (
    addr_width_b => 8,
    clocking_mode => "common_clock",
    data_width_b => 18,
    latency => 1,
    mem_init_file => "xpm_d42629_vivado.mem",
    mem_size => 4608,
    mem_type => "block",
    read_reset_a => "0",
    read_reset_b => "0",
    width => 18,
    width_addr => 8,
    write_mode_a => "read_first",
    write_mode_b => "read_first"
  )
  port map (
    ena => "1",
    enb => "1",
    rsta => "0",
    rstb => "0",
    addra => ram_dphi_addr_op_net,
    dina => constant3_op_net,
    wea => constant_op_net,
    addrb => delay38_q_net,
    dinb => delay44_q_net,
    web => delay49_q_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dpram_init_im_even_4_douta_net,
    doutb => dpram_init_im_even_4_doutb_net
  );
  dpram_init_re_even_4 : entity xil_defaultlib.psb3_0_xltdpram 
  generic map (
    addr_width_b => 8,
    clocking_mode => "common_clock",
    data_width_b => 18,
    latency => 1,
    mem_init_file => "xpm_3895d5_vivado.mem",
    mem_size => 4608,
    mem_type => "block",
    read_reset_a => "0",
    read_reset_b => "0",
    width => 18,
    width_addr => 8,
    write_mode_a => "read_first",
    write_mode_b => "read_first"
  )
  port map (
    ena => "1",
    enb => "1",
    rsta => "0",
    rstb => "0",
    addra => ram_dphi_addr_op_net,
    dina => constant7_op_net,
    wea => constant1_op_net,
    addrb => delay38_q_net,
    dinb => delay35_q_net,
    web => delay49_q_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dpram_init_re_even_4_douta_net,
    doutb => dpram_init_re_even_4_doutb_net
  );
  delay16 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 253,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => constant6_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay16_q_net
  );
  fifo4 : entity xil_defaultlib.psb3_0_xlfifogen_u 
  generic map (
    core_name0 => "psb3_0_fifo_generator_i1",
    data_count_width => 10,
    data_width => 16,
    extra_registers => 1,
    has_ae => 0,
    has_af => 0,
    has_rst => false,
    ignore_din_for_gcd => false,
    percent_full_width => 1
  )
  port map (
    en => '1',
    rst => '0',
    din => addsub_s_net,
    we => constant6_op_net(0),
    re => delay16_q_net(0),
    clk => clk_net,
    ce => ce_net,
    we_ce => ce_net,
    re_ce => ce_net,
    dout => fifo4_dout_net,
    empty => fifo4_empty_net,
    full => fifo4_full_net
  );
  reinterpret2 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => fifo4_dout_net,
    output_port => reinterpret2_output_port_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Baseband_odd_1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_baseband_odd_1 is
  port (
    tvalid : in std_logic_vector( 1-1 downto 0 );
    addr_r : in std_logic_vector( 8-1 downto 0 );
    addr_w : in std_logic_vector( 8-1 downto 0 );
    init_im_odd : in std_logic_vector( 18-1 downto 0 );
    init_re_odd : in std_logic_vector( 18-1 downto 0 );
    dphi_odd : in std_logic_vector( 16-1 downto 0 );
    we : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    out_im : out std_logic_vector( 16-1 downto 0 );
    out_re : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_baseband_odd_1;
architecture structural of psb3_0_baseband_odd_1 is 
  signal cordic_6_0_odd_1_m_axis_dout_tdata_imag_net : std_logic_vector( 16-1 downto 0 );
  signal cordic_6_0_odd_1_m_axis_dout_tdata_real_net : std_logic_vector( 16-1 downto 0 );
  signal delay37_q_net : std_logic_vector( 16-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay44_q_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal dpram_dphi_odd_1_douta_net : std_logic_vector( 16-1 downto 0 );
  signal cordic_6_0_odd_1_m_axis_dout_tvalid_net : std_logic;
  signal delay14_q_net : std_logic_vector( 1-1 downto 0 );
  signal ram_dphi_addr_op_net : std_logic_vector( 8-1 downto 0 );
  signal delay35_q_net : std_logic_vector( 18-1 downto 0 );
  signal fifo1_dout_net : std_logic_vector( 16-1 downto 0 );
  signal delay38_q_net : std_logic_vector( 8-1 downto 0 );
  signal ce_net : std_logic;
  signal addsub1_s_net : std_logic_vector( 16-1 downto 0 );
  signal dpram_init_im_odd_1_douta_net : std_logic_vector( 18-1 downto 0 );
  signal dpram_init_re_odd_1_douta_net : std_logic_vector( 18-1 downto 0 );
  signal convert1_dout_net : std_logic_vector( 18-1 downto 0 );
  signal constant10_op_net : std_logic_vector( 18-1 downto 0 );
  signal constant5_op_net : std_logic_vector( 1-1 downto 0 );
  signal dpram_dphi_odd_1_doutb_net : std_logic_vector( 16-1 downto 0 );
  signal constant12_op_net : std_logic_vector( 18-1 downto 0 );
  signal constant13_op_net : std_logic_vector( 16-1 downto 0 );
  signal constant4_op_net : std_logic_vector( 1-1 downto 0 );
  signal constant11_op_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal constant9_op_net : std_logic_vector( 1-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 1-1 downto 0 );
  signal dpram_init_im_odd_1_doutb_net : std_logic_vector( 18-1 downto 0 );
  signal dpram_init_re_odd_1_doutb_net : std_logic_vector( 18-1 downto 0 );
  signal fifo1_full_net : std_logic;
  signal fifo1_empty_net : std_logic;
begin
  out_im <= cordic_6_0_odd_1_m_axis_dout_tdata_imag_net;
  out_re <= cordic_6_0_odd_1_m_axis_dout_tdata_real_net;
  delay14_q_net <= tvalid;
  ram_dphi_addr_op_net <= addr_r;
  delay38_q_net <= addr_w;
  delay44_q_net <= init_im_odd;
  delay35_q_net <= init_re_odd;
  delay37_q_net <= dphi_odd;
  delay6_q_net <= we;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub1 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 16,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 17,
    core_name0 => "psb3_0_c_addsub_v12_0_i0",
    extra_registers => 1,
    full_s_arith => 1,
    full_s_width => 17,
    latency => 2,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => dpram_dphi_odd_1_douta_net,
    b => fifo1_dout_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  cordic_6_0_odd_1 : entity xil_defaultlib.xlcordic_5a76bbdd6458ef1eb96e9ff32fab9279 
  port map (
    s_axis_cartesian_tvalid => delay14_q_net(0),
    s_axis_cartesian_tdata_imag => dpram_init_im_odd_1_douta_net,
    s_axis_cartesian_tdata_real => dpram_init_re_odd_1_douta_net,
    s_axis_phase_tvalid => delay14_q_net(0),
    s_axis_phase_tdata_phase => convert1_dout_net,
    clk => clk_net,
    ce => ce_net,
    m_axis_dout_tvalid => cordic_6_0_odd_1_m_axis_dout_tvalid_net,
    m_axis_dout_tdata_imag => cordic_6_0_odd_1_m_axis_dout_tdata_imag_net,
    m_axis_dout_tdata_real => cordic_6_0_odd_1_m_axis_dout_tdata_real_net
  );
  constant10 : entity xil_defaultlib.sysgen_constant_ac4aa5284f 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant10_op_net
  );
  constant11 : entity xil_defaultlib.sysgen_constant_71e89d757c 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant11_op_net
  );
  constant12 : entity xil_defaultlib.sysgen_constant_ac4aa5284f 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant12_op_net
  );
  constant13 : entity xil_defaultlib.sysgen_constant_eb74b92b90 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant13_op_net
  );
  constant4 : entity xil_defaultlib.sysgen_constant_de9059c03f 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant4_op_net
  );
  constant5 : entity xil_defaultlib.sysgen_constant_de9059c03f 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant5_op_net
  );
  constant9 : entity xil_defaultlib.sysgen_constant_de9059c03f 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant9_op_net
  );
  convert1 : entity xil_defaultlib.psb3_0_xlconvert 
  generic map (
    bool_conversion => 0,
    din_arith => 2,
    din_bin_pt => 15,
    din_width => 16,
    dout_arith => 2,
    dout_bin_pt => 15,
    dout_width => 18,
    latency => 0,
    overflow => xlWrap,
    quantization => xlTruncate
  )
  port map (
    clr => '0',
    en => "1",
    din => reinterpret1_output_port_net,
    clk => clk_net,
    ce => ce_net,
    dout => convert1_dout_net
  );
  dpram_dphi_odd_1 : entity xil_defaultlib.psb3_0_xltdpram 
  generic map (
    addr_width_b => 8,
    clocking_mode => "common_clock",
    data_width_b => 16,
    latency => 1,
    mem_init_file => "xpm_95ed83_vivado.mem",
    mem_size => 4096,
    mem_type => "block",
    read_reset_a => "0",
    read_reset_b => "0",
    width => 16,
    width_addr => 8,
    write_mode_a => "read_first",
    write_mode_b => "read_first"
  )
  port map (
    ena => "1",
    enb => "1",
    rsta => "0",
    rstb => "0",
    addra => ram_dphi_addr_op_net,
    dina => constant13_op_net,
    wea => constant9_op_net,
    addrb => delay38_q_net,
    dinb => delay37_q_net,
    web => delay6_q_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dpram_dphi_odd_1_douta_net,
    doutb => dpram_dphi_odd_1_doutb_net
  );
  dpram_init_im_odd_1 : entity xil_defaultlib.psb3_0_xltdpram 
  generic map (
    addr_width_b => 8,
    clocking_mode => "common_clock",
    data_width_b => 18,
    latency => 1,
    mem_init_file => "xpm_d15418_vivado.mem",
    mem_size => 4608,
    mem_type => "block",
    read_reset_a => "0",
    read_reset_b => "0",
    width => 18,
    width_addr => 8,
    write_mode_a => "read_first",
    write_mode_b => "read_first"
  )
  port map (
    ena => "1",
    enb => "1",
    rsta => "0",
    rstb => "0",
    addra => ram_dphi_addr_op_net,
    dina => constant10_op_net,
    wea => constant4_op_net,
    addrb => delay38_q_net,
    dinb => delay44_q_net,
    web => delay6_q_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dpram_init_im_odd_1_douta_net,
    doutb => dpram_init_im_odd_1_doutb_net
  );
  dpram_init_re_odd_1 : entity xil_defaultlib.psb3_0_xltdpram 
  generic map (
    addr_width_b => 8,
    clocking_mode => "common_clock",
    data_width_b => 18,
    latency => 1,
    mem_init_file => "xpm_2f56aa_vivado.mem",
    mem_size => 4608,
    mem_type => "block",
    read_reset_a => "0",
    read_reset_b => "0",
    width => 18,
    width_addr => 8,
    write_mode_a => "read_first",
    write_mode_b => "read_first"
  )
  port map (
    ena => "1",
    enb => "1",
    rsta => "0",
    rstb => "0",
    addra => ram_dphi_addr_op_net,
    dina => constant12_op_net,
    wea => constant5_op_net,
    addrb => delay38_q_net,
    dinb => delay35_q_net,
    web => delay6_q_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dpram_init_re_odd_1_douta_net,
    doutb => dpram_init_re_odd_1_doutb_net
  );
  delay8 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 253,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => constant11_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay8_q_net
  );
  fifo1 : entity xil_defaultlib.psb3_0_xlfifogen_u 
  generic map (
    core_name0 => "psb3_0_fifo_generator_i1",
    data_count_width => 10,
    data_width => 16,
    extra_registers => 1,
    has_ae => 0,
    has_af => 0,
    has_rst => false,
    ignore_din_for_gcd => false,
    percent_full_width => 1
  )
  port map (
    en => '1',
    rst => '0',
    din => addsub1_s_net,
    we => constant11_op_net(0),
    re => delay8_q_net(0),
    clk => clk_net,
    ce => ce_net,
    we_ce => ce_net,
    re_ce => ce_net,
    dout => fifo1_dout_net,
    empty => fifo1_empty_net,
    full => fifo1_full_net
  );
  reinterpret1 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => fifo1_dout_net,
    output_port => reinterpret1_output_port_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Baseband_odd_2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_baseband_odd_2 is
  port (
    tvalid : in std_logic_vector( 1-1 downto 0 );
    addr_r : in std_logic_vector( 8-1 downto 0 );
    addr_w : in std_logic_vector( 8-1 downto 0 );
    init_im_odd_2 : in std_logic_vector( 18-1 downto 0 );
    init_re_odd_2 : in std_logic_vector( 18-1 downto 0 );
    dphi_odd_2 : in std_logic_vector( 16-1 downto 0 );
    we : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    out_im : out std_logic_vector( 16-1 downto 0 );
    out_re : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_baseband_odd_2;
architecture structural of psb3_0_baseband_odd_2 is 
  signal addsub1_s_net : std_logic_vector( 16-1 downto 0 );
  signal delay26_q_net : std_logic_vector( 1-1 downto 0 );
  signal dpram_dphi_odd_2_douta_net : std_logic_vector( 16-1 downto 0 );
  signal delay35_q_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal ram_dphi_addr_op_net : std_logic_vector( 8-1 downto 0 );
  signal delay38_q_net : std_logic_vector( 8-1 downto 0 );
  signal delay14_q_net : std_logic_vector( 1-1 downto 0 );
  signal fifo1_dout_net : std_logic_vector( 16-1 downto 0 );
  signal delay44_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay37_q_net : std_logic_vector( 16-1 downto 0 );
  signal clk_net : std_logic;
  signal cordic_6_0_odd_2_m_axis_dout_tdata_imag_net : std_logic_vector( 16-1 downto 0 );
  signal cordic_6_0_odd_2_m_axis_dout_tdata_real_net : std_logic_vector( 16-1 downto 0 );
  signal constant10_op_net : std_logic_vector( 18-1 downto 0 );
  signal constant11_op_net : std_logic_vector( 1-1 downto 0 );
  signal dpram_init_im_odd_2_douta_net : std_logic_vector( 18-1 downto 0 );
  signal constant13_op_net : std_logic_vector( 16-1 downto 0 );
  signal dpram_init_re_odd_2_douta_net : std_logic_vector( 18-1 downto 0 );
  signal convert1_dout_net : std_logic_vector( 18-1 downto 0 );
  signal constant4_op_net : std_logic_vector( 1-1 downto 0 );
  signal constant12_op_net : std_logic_vector( 18-1 downto 0 );
  signal constant5_op_net : std_logic_vector( 1-1 downto 0 );
  signal constant9_op_net : std_logic_vector( 1-1 downto 0 );
  signal cordic_6_0_odd_2_m_axis_dout_tvalid_net : std_logic;
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal dpram_init_im_odd_2_doutb_net : std_logic_vector( 18-1 downto 0 );
  signal dpram_init_re_odd_2_doutb_net : std_logic_vector( 18-1 downto 0 );
  signal dpram_dphi_odd_2_doutb_net : std_logic_vector( 16-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 1-1 downto 0 );
  signal fifo1_full_net : std_logic;
  signal fifo1_empty_net : std_logic;
begin
  out_im <= cordic_6_0_odd_2_m_axis_dout_tdata_imag_net;
  out_re <= cordic_6_0_odd_2_m_axis_dout_tdata_real_net;
  delay14_q_net <= tvalid;
  ram_dphi_addr_op_net <= addr_r;
  delay38_q_net <= addr_w;
  delay44_q_net <= init_im_odd_2;
  delay35_q_net <= init_re_odd_2;
  delay37_q_net <= dphi_odd_2;
  delay26_q_net <= we;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub1 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 16,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 17,
    core_name0 => "psb3_0_c_addsub_v12_0_i0",
    extra_registers => 1,
    full_s_arith => 1,
    full_s_width => 17,
    latency => 2,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => dpram_dphi_odd_2_douta_net,
    b => fifo1_dout_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  cordic_6_0_odd_2 : entity xil_defaultlib.xlcordic_5a76bbdd6458ef1eb96e9ff32fab9279 
  port map (
    s_axis_cartesian_tvalid => delay14_q_net(0),
    s_axis_cartesian_tdata_imag => dpram_init_im_odd_2_douta_net,
    s_axis_cartesian_tdata_real => dpram_init_re_odd_2_douta_net,
    s_axis_phase_tvalid => delay14_q_net(0),
    s_axis_phase_tdata_phase => convert1_dout_net,
    clk => clk_net,
    ce => ce_net,
    m_axis_dout_tvalid => cordic_6_0_odd_2_m_axis_dout_tvalid_net,
    m_axis_dout_tdata_imag => cordic_6_0_odd_2_m_axis_dout_tdata_imag_net,
    m_axis_dout_tdata_real => cordic_6_0_odd_2_m_axis_dout_tdata_real_net
  );
  constant10 : entity xil_defaultlib.sysgen_constant_ac4aa5284f 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant10_op_net
  );
  constant11 : entity xil_defaultlib.sysgen_constant_71e89d757c 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant11_op_net
  );
  constant12 : entity xil_defaultlib.sysgen_constant_ac4aa5284f 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant12_op_net
  );
  constant13 : entity xil_defaultlib.sysgen_constant_eb74b92b90 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant13_op_net
  );
  constant4 : entity xil_defaultlib.sysgen_constant_de9059c03f 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant4_op_net
  );
  constant5 : entity xil_defaultlib.sysgen_constant_de9059c03f 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant5_op_net
  );
  constant9 : entity xil_defaultlib.sysgen_constant_de9059c03f 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant9_op_net
  );
  convert1 : entity xil_defaultlib.psb3_0_xlconvert 
  generic map (
    bool_conversion => 0,
    din_arith => 2,
    din_bin_pt => 15,
    din_width => 16,
    dout_arith => 2,
    dout_bin_pt => 15,
    dout_width => 18,
    latency => 0,
    overflow => xlWrap,
    quantization => xlTruncate
  )
  port map (
    clr => '0',
    en => "1",
    din => reinterpret1_output_port_net,
    clk => clk_net,
    ce => ce_net,
    dout => convert1_dout_net
  );
  dpram_dphi_odd_2 : entity xil_defaultlib.psb3_0_xltdpram 
  generic map (
    addr_width_b => 8,
    clocking_mode => "common_clock",
    data_width_b => 16,
    latency => 1,
    mem_init_file => "xpm_c4fac8_vivado.mem",
    mem_size => 4096,
    mem_type => "block",
    read_reset_a => "0",
    read_reset_b => "0",
    width => 16,
    width_addr => 8,
    write_mode_a => "read_first",
    write_mode_b => "read_first"
  )
  port map (
    ena => "1",
    enb => "1",
    rsta => "0",
    rstb => "0",
    addra => ram_dphi_addr_op_net,
    dina => constant13_op_net,
    wea => constant9_op_net,
    addrb => delay38_q_net,
    dinb => delay37_q_net,
    web => delay26_q_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dpram_dphi_odd_2_douta_net,
    doutb => dpram_dphi_odd_2_doutb_net
  );
  dpram_init_im_odd_2 : entity xil_defaultlib.psb3_0_xltdpram 
  generic map (
    addr_width_b => 8,
    clocking_mode => "common_clock",
    data_width_b => 18,
    latency => 1,
    mem_init_file => "xpm_8b0ba2_vivado.mem",
    mem_size => 4608,
    mem_type => "block",
    read_reset_a => "0",
    read_reset_b => "0",
    width => 18,
    width_addr => 8,
    write_mode_a => "read_first",
    write_mode_b => "read_first"
  )
  port map (
    ena => "1",
    enb => "1",
    rsta => "0",
    rstb => "0",
    addra => ram_dphi_addr_op_net,
    dina => constant10_op_net,
    wea => constant4_op_net,
    addrb => delay38_q_net,
    dinb => delay44_q_net,
    web => delay26_q_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dpram_init_im_odd_2_douta_net,
    doutb => dpram_init_im_odd_2_doutb_net
  );
  dpram_init_re_odd_2 : entity xil_defaultlib.psb3_0_xltdpram 
  generic map (
    addr_width_b => 8,
    clocking_mode => "common_clock",
    data_width_b => 18,
    latency => 1,
    mem_init_file => "xpm_6cb1ed_vivado.mem",
    mem_size => 4608,
    mem_type => "block",
    read_reset_a => "0",
    read_reset_b => "0",
    width => 18,
    width_addr => 8,
    write_mode_a => "read_first",
    write_mode_b => "read_first"
  )
  port map (
    ena => "1",
    enb => "1",
    rsta => "0",
    rstb => "0",
    addra => ram_dphi_addr_op_net,
    dina => constant12_op_net,
    wea => constant5_op_net,
    addrb => delay38_q_net,
    dinb => delay35_q_net,
    web => delay26_q_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dpram_init_re_odd_2_douta_net,
    doutb => dpram_init_re_odd_2_doutb_net
  );
  delay8 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 253,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => constant11_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay8_q_net
  );
  fifo1 : entity xil_defaultlib.psb3_0_xlfifogen_u 
  generic map (
    core_name0 => "psb3_0_fifo_generator_i1",
    data_count_width => 10,
    data_width => 16,
    extra_registers => 1,
    has_ae => 0,
    has_af => 0,
    has_rst => false,
    ignore_din_for_gcd => false,
    percent_full_width => 1
  )
  port map (
    en => '1',
    rst => '0',
    din => addsub1_s_net,
    we => constant11_op_net(0),
    re => delay8_q_net(0),
    clk => clk_net,
    ce => ce_net,
    we_ce => ce_net,
    re_ce => ce_net,
    dout => fifo1_dout_net,
    empty => fifo1_empty_net,
    full => fifo1_full_net
  );
  reinterpret1 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => fifo1_dout_net,
    output_port => reinterpret1_output_port_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Baseband_odd_3
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_baseband_odd_3 is
  port (
    tvalid : in std_logic_vector( 1-1 downto 0 );
    addr_r : in std_logic_vector( 8-1 downto 0 );
    addr_w : in std_logic_vector( 8-1 downto 0 );
    init_im_odd : in std_logic_vector( 18-1 downto 0 );
    init_re_odd : in std_logic_vector( 18-1 downto 0 );
    dphi_odd : in std_logic_vector( 16-1 downto 0 );
    we : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    out_im : out std_logic_vector( 16-1 downto 0 );
    out_re : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_baseband_odd_3;
architecture structural of psb3_0_baseband_odd_3 is 
  signal delay35_q_net : std_logic_vector( 18-1 downto 0 );
  signal cordic_6_0_odd_1_m_axis_dout_tdata_imag_net : std_logic_vector( 16-1 downto 0 );
  signal delay44_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay37_q_net : std_logic_vector( 16-1 downto 0 );
  signal delay14_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay38_q_net : std_logic_vector( 8-1 downto 0 );
  signal clk_net : std_logic;
  signal cordic_6_0_odd_1_m_axis_dout_tdata_real_net : std_logic_vector( 16-1 downto 0 );
  signal ram_dphi_addr_op_net : std_logic_vector( 8-1 downto 0 );
  signal delay48_q_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal addsub1_s_net : std_logic_vector( 16-1 downto 0 );
  signal dpram_init_re_odd_3_douta_net : std_logic_vector( 18-1 downto 0 );
  signal constant12_op_net : std_logic_vector( 18-1 downto 0 );
  signal dpram_dphi_odd_3_douta_net : std_logic_vector( 16-1 downto 0 );
  signal convert1_dout_net : std_logic_vector( 18-1 downto 0 );
  signal dpram_init_im_odd_3_douta_net : std_logic_vector( 18-1 downto 0 );
  signal constant13_op_net : std_logic_vector( 16-1 downto 0 );
  signal constant10_op_net : std_logic_vector( 18-1 downto 0 );
  signal constant5_op_net : std_logic_vector( 1-1 downto 0 );
  signal constant4_op_net : std_logic_vector( 1-1 downto 0 );
  signal fifo1_dout_net : std_logic_vector( 16-1 downto 0 );
  signal constant11_op_net : std_logic_vector( 1-1 downto 0 );
  signal cordic_6_0_odd_1_m_axis_dout_tvalid_net : std_logic;
  signal dpram_dphi_odd_3_doutb_net : std_logic_vector( 16-1 downto 0 );
  signal constant9_op_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal dpram_init_im_odd_3_doutb_net : std_logic_vector( 18-1 downto 0 );
  signal dpram_init_re_odd_3_doutb_net : std_logic_vector( 18-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 1-1 downto 0 );
  signal fifo1_full_net : std_logic;
  signal fifo1_empty_net : std_logic;
begin
  out_im <= cordic_6_0_odd_1_m_axis_dout_tdata_imag_net;
  out_re <= cordic_6_0_odd_1_m_axis_dout_tdata_real_net;
  delay14_q_net <= tvalid;
  ram_dphi_addr_op_net <= addr_r;
  delay38_q_net <= addr_w;
  delay44_q_net <= init_im_odd;
  delay35_q_net <= init_re_odd;
  delay37_q_net <= dphi_odd;
  delay48_q_net <= we;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub1 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 16,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 17,
    core_name0 => "psb3_0_c_addsub_v12_0_i0",
    extra_registers => 1,
    full_s_arith => 1,
    full_s_width => 17,
    latency => 2,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => dpram_dphi_odd_3_douta_net,
    b => fifo1_dout_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  cordic_6_0_odd_1 : entity xil_defaultlib.xlcordic_5a76bbdd6458ef1eb96e9ff32fab9279 
  port map (
    s_axis_cartesian_tvalid => delay14_q_net(0),
    s_axis_cartesian_tdata_imag => dpram_init_im_odd_3_douta_net,
    s_axis_cartesian_tdata_real => dpram_init_re_odd_3_douta_net,
    s_axis_phase_tvalid => delay14_q_net(0),
    s_axis_phase_tdata_phase => convert1_dout_net,
    clk => clk_net,
    ce => ce_net,
    m_axis_dout_tvalid => cordic_6_0_odd_1_m_axis_dout_tvalid_net,
    m_axis_dout_tdata_imag => cordic_6_0_odd_1_m_axis_dout_tdata_imag_net,
    m_axis_dout_tdata_real => cordic_6_0_odd_1_m_axis_dout_tdata_real_net
  );
  constant10 : entity xil_defaultlib.sysgen_constant_ac4aa5284f 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant10_op_net
  );
  constant11 : entity xil_defaultlib.sysgen_constant_71e89d757c 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant11_op_net
  );
  constant12 : entity xil_defaultlib.sysgen_constant_ac4aa5284f 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant12_op_net
  );
  constant13 : entity xil_defaultlib.sysgen_constant_eb74b92b90 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant13_op_net
  );
  constant4 : entity xil_defaultlib.sysgen_constant_de9059c03f 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant4_op_net
  );
  constant5 : entity xil_defaultlib.sysgen_constant_de9059c03f 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant5_op_net
  );
  constant9 : entity xil_defaultlib.sysgen_constant_de9059c03f 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant9_op_net
  );
  convert1 : entity xil_defaultlib.psb3_0_xlconvert 
  generic map (
    bool_conversion => 0,
    din_arith => 2,
    din_bin_pt => 15,
    din_width => 16,
    dout_arith => 2,
    dout_bin_pt => 15,
    dout_width => 18,
    latency => 0,
    overflow => xlWrap,
    quantization => xlTruncate
  )
  port map (
    clr => '0',
    en => "1",
    din => reinterpret1_output_port_net,
    clk => clk_net,
    ce => ce_net,
    dout => convert1_dout_net
  );
  dpram_dphi_odd_3 : entity xil_defaultlib.psb3_0_xltdpram 
  generic map (
    addr_width_b => 8,
    clocking_mode => "common_clock",
    data_width_b => 16,
    latency => 1,
    mem_init_file => "xpm_8ca7ae_vivado.mem",
    mem_size => 4096,
    mem_type => "block",
    read_reset_a => "0",
    read_reset_b => "0",
    width => 16,
    width_addr => 8,
    write_mode_a => "read_first",
    write_mode_b => "read_first"
  )
  port map (
    ena => "1",
    enb => "1",
    rsta => "0",
    rstb => "0",
    addra => ram_dphi_addr_op_net,
    dina => constant13_op_net,
    wea => constant9_op_net,
    addrb => delay38_q_net,
    dinb => delay37_q_net,
    web => delay48_q_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dpram_dphi_odd_3_douta_net,
    doutb => dpram_dphi_odd_3_doutb_net
  );
  dpram_init_im_odd_3 : entity xil_defaultlib.psb3_0_xltdpram 
  generic map (
    addr_width_b => 8,
    clocking_mode => "common_clock",
    data_width_b => 18,
    latency => 1,
    mem_init_file => "xpm_53a103_vivado.mem",
    mem_size => 4608,
    mem_type => "block",
    read_reset_a => "0",
    read_reset_b => "0",
    width => 18,
    width_addr => 8,
    write_mode_a => "read_first",
    write_mode_b => "read_first"
  )
  port map (
    ena => "1",
    enb => "1",
    rsta => "0",
    rstb => "0",
    addra => ram_dphi_addr_op_net,
    dina => constant10_op_net,
    wea => constant4_op_net,
    addrb => delay38_q_net,
    dinb => delay44_q_net,
    web => delay48_q_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dpram_init_im_odd_3_douta_net,
    doutb => dpram_init_im_odd_3_doutb_net
  );
  dpram_init_re_odd_3 : entity xil_defaultlib.psb3_0_xltdpram 
  generic map (
    addr_width_b => 8,
    clocking_mode => "common_clock",
    data_width_b => 18,
    latency => 1,
    mem_init_file => "xpm_196cb0_vivado.mem",
    mem_size => 4608,
    mem_type => "block",
    read_reset_a => "0",
    read_reset_b => "0",
    width => 18,
    width_addr => 8,
    write_mode_a => "read_first",
    write_mode_b => "read_first"
  )
  port map (
    ena => "1",
    enb => "1",
    rsta => "0",
    rstb => "0",
    addra => ram_dphi_addr_op_net,
    dina => constant12_op_net,
    wea => constant5_op_net,
    addrb => delay38_q_net,
    dinb => delay35_q_net,
    web => delay48_q_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dpram_init_re_odd_3_douta_net,
    doutb => dpram_init_re_odd_3_doutb_net
  );
  delay8 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 253,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => constant11_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay8_q_net
  );
  fifo1 : entity xil_defaultlib.psb3_0_xlfifogen_u 
  generic map (
    core_name0 => "psb3_0_fifo_generator_i1",
    data_count_width => 10,
    data_width => 16,
    extra_registers => 1,
    has_ae => 0,
    has_af => 0,
    has_rst => false,
    ignore_din_for_gcd => false,
    percent_full_width => 1
  )
  port map (
    en => '1',
    rst => '0',
    din => addsub1_s_net,
    we => constant11_op_net(0),
    re => delay8_q_net(0),
    clk => clk_net,
    ce => ce_net,
    we_ce => ce_net,
    re_ce => ce_net,
    dout => fifo1_dout_net,
    empty => fifo1_empty_net,
    full => fifo1_full_net
  );
  reinterpret1 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => fifo1_dout_net,
    output_port => reinterpret1_output_port_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Baseband_odd_4
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_baseband_odd_4 is
  port (
    tvalid : in std_logic_vector( 1-1 downto 0 );
    addr_r : in std_logic_vector( 8-1 downto 0 );
    addr_w : in std_logic_vector( 8-1 downto 0 );
    init_im_odd_2 : in std_logic_vector( 18-1 downto 0 );
    init_re_odd_2 : in std_logic_vector( 18-1 downto 0 );
    dphi_odd_2 : in std_logic_vector( 16-1 downto 0 );
    we : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    out_im : out std_logic_vector( 16-1 downto 0 );
    out_re : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_baseband_odd_4;
architecture structural of psb3_0_baseband_odd_4 is 
  signal ram_dphi_addr_op_net : std_logic_vector( 8-1 downto 0 );
  signal delay44_q_net : std_logic_vector( 18-1 downto 0 );
  signal cordic_6_0_odd_2_m_axis_dout_tdata_real_net : std_logic_vector( 16-1 downto 0 );
  signal delay14_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay38_q_net : std_logic_vector( 8-1 downto 0 );
  signal delay35_q_net : std_logic_vector( 18-1 downto 0 );
  signal cordic_6_0_odd_2_m_axis_dout_tdata_imag_net : std_logic_vector( 16-1 downto 0 );
  signal delay37_q_net : std_logic_vector( 16-1 downto 0 );
  signal delay43_q_net : std_logic_vector( 1-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 16-1 downto 0 );
  signal ce_net : std_logic;
  signal clk_net : std_logic;
  signal dpram_dphi_odd_4_douta_net : std_logic_vector( 16-1 downto 0 );
  signal fifo1_dout_net : std_logic_vector( 16-1 downto 0 );
  signal dpram_init_re_odd_4_douta_net : std_logic_vector( 18-1 downto 0 );
  signal convert1_dout_net : std_logic_vector( 18-1 downto 0 );
  signal dpram_init_im_odd_4_douta_net : std_logic_vector( 18-1 downto 0 );
  signal cordic_6_0_odd_2_m_axis_dout_tvalid_net : std_logic;
  signal constant10_op_net : std_logic_vector( 18-1 downto 0 );
  signal constant11_op_net : std_logic_vector( 1-1 downto 0 );
  signal constant12_op_net : std_logic_vector( 18-1 downto 0 );
  signal constant4_op_net : std_logic_vector( 1-1 downto 0 );
  signal constant13_op_net : std_logic_vector( 16-1 downto 0 );
  signal constant9_op_net : std_logic_vector( 1-1 downto 0 );
  signal constant5_op_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal dpram_dphi_odd_4_doutb_net : std_logic_vector( 16-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 1-1 downto 0 );
  signal dpram_init_re_odd_4_doutb_net : std_logic_vector( 18-1 downto 0 );
  signal dpram_init_im_odd_4_doutb_net : std_logic_vector( 18-1 downto 0 );
  signal fifo1_empty_net : std_logic;
  signal fifo1_full_net : std_logic;
begin
  out_im <= cordic_6_0_odd_2_m_axis_dout_tdata_imag_net;
  out_re <= cordic_6_0_odd_2_m_axis_dout_tdata_real_net;
  delay14_q_net <= tvalid;
  ram_dphi_addr_op_net <= addr_r;
  delay38_q_net <= addr_w;
  delay44_q_net <= init_im_odd_2;
  delay35_q_net <= init_re_odd_2;
  delay37_q_net <= dphi_odd_2;
  delay43_q_net <= we;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub1 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 16,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 17,
    core_name0 => "psb3_0_c_addsub_v12_0_i0",
    extra_registers => 1,
    full_s_arith => 1,
    full_s_width => 17,
    latency => 2,
    overflow => 1,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => dpram_dphi_odd_4_douta_net,
    b => fifo1_dout_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  cordic_6_0_odd_2 : entity xil_defaultlib.xlcordic_5a76bbdd6458ef1eb96e9ff32fab9279 
  port map (
    s_axis_cartesian_tvalid => delay14_q_net(0),
    s_axis_cartesian_tdata_imag => dpram_init_im_odd_4_douta_net,
    s_axis_cartesian_tdata_real => dpram_init_re_odd_4_douta_net,
    s_axis_phase_tvalid => delay14_q_net(0),
    s_axis_phase_tdata_phase => convert1_dout_net,
    clk => clk_net,
    ce => ce_net,
    m_axis_dout_tvalid => cordic_6_0_odd_2_m_axis_dout_tvalid_net,
    m_axis_dout_tdata_imag => cordic_6_0_odd_2_m_axis_dout_tdata_imag_net,
    m_axis_dout_tdata_real => cordic_6_0_odd_2_m_axis_dout_tdata_real_net
  );
  constant10 : entity xil_defaultlib.sysgen_constant_ac4aa5284f 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant10_op_net
  );
  constant11 : entity xil_defaultlib.sysgen_constant_71e89d757c 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant11_op_net
  );
  constant12 : entity xil_defaultlib.sysgen_constant_ac4aa5284f 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant12_op_net
  );
  constant13 : entity xil_defaultlib.sysgen_constant_eb74b92b90 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant13_op_net
  );
  constant4 : entity xil_defaultlib.sysgen_constant_de9059c03f 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant4_op_net
  );
  constant5 : entity xil_defaultlib.sysgen_constant_de9059c03f 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant5_op_net
  );
  constant9 : entity xil_defaultlib.sysgen_constant_de9059c03f 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant9_op_net
  );
  convert1 : entity xil_defaultlib.psb3_0_xlconvert 
  generic map (
    bool_conversion => 0,
    din_arith => 2,
    din_bin_pt => 15,
    din_width => 16,
    dout_arith => 2,
    dout_bin_pt => 15,
    dout_width => 18,
    latency => 0,
    overflow => xlWrap,
    quantization => xlTruncate
  )
  port map (
    clr => '0',
    en => "1",
    din => reinterpret1_output_port_net,
    clk => clk_net,
    ce => ce_net,
    dout => convert1_dout_net
  );
  dpram_dphi_odd_4 : entity xil_defaultlib.psb3_0_xltdpram 
  generic map (
    addr_width_b => 8,
    clocking_mode => "common_clock",
    data_width_b => 16,
    latency => 1,
    mem_init_file => "xpm_d23bbc_vivado.mem",
    mem_size => 4096,
    mem_type => "block",
    read_reset_a => "0",
    read_reset_b => "0",
    width => 16,
    width_addr => 8,
    write_mode_a => "read_first",
    write_mode_b => "read_first"
  )
  port map (
    ena => "1",
    enb => "1",
    rsta => "0",
    rstb => "0",
    addra => ram_dphi_addr_op_net,
    dina => constant13_op_net,
    wea => constant9_op_net,
    addrb => delay38_q_net,
    dinb => delay37_q_net,
    web => delay43_q_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dpram_dphi_odd_4_douta_net,
    doutb => dpram_dphi_odd_4_doutb_net
  );
  dpram_init_im_odd_4 : entity xil_defaultlib.psb3_0_xltdpram 
  generic map (
    addr_width_b => 8,
    clocking_mode => "common_clock",
    data_width_b => 18,
    latency => 1,
    mem_init_file => "xpm_fb9180_vivado.mem",
    mem_size => 4608,
    mem_type => "block",
    read_reset_a => "0",
    read_reset_b => "0",
    width => 18,
    width_addr => 8,
    write_mode_a => "read_first",
    write_mode_b => "read_first"
  )
  port map (
    ena => "1",
    enb => "1",
    rsta => "0",
    rstb => "0",
    addra => ram_dphi_addr_op_net,
    dina => constant10_op_net,
    wea => constant4_op_net,
    addrb => delay38_q_net,
    dinb => delay44_q_net,
    web => delay43_q_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dpram_init_im_odd_4_douta_net,
    doutb => dpram_init_im_odd_4_doutb_net
  );
  dpram_init_re_odd_4 : entity xil_defaultlib.psb3_0_xltdpram 
  generic map (
    addr_width_b => 8,
    clocking_mode => "common_clock",
    data_width_b => 18,
    latency => 1,
    mem_init_file => "xpm_db9fae_vivado.mem",
    mem_size => 4608,
    mem_type => "block",
    read_reset_a => "0",
    read_reset_b => "0",
    width => 18,
    width_addr => 8,
    write_mode_a => "read_first",
    write_mode_b => "read_first"
  )
  port map (
    ena => "1",
    enb => "1",
    rsta => "0",
    rstb => "0",
    addra => ram_dphi_addr_op_net,
    dina => constant12_op_net,
    wea => constant5_op_net,
    addrb => delay38_q_net,
    dinb => delay35_q_net,
    web => delay43_q_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dpram_init_re_odd_4_douta_net,
    doutb => dpram_init_re_odd_4_doutb_net
  );
  delay8 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 253,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => constant11_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay8_q_net
  );
  fifo1 : entity xil_defaultlib.psb3_0_xlfifogen_u 
  generic map (
    core_name0 => "psb3_0_fifo_generator_i1",
    data_count_width => 10,
    data_width => 16,
    extra_registers => 1,
    has_ae => 0,
    has_af => 0,
    has_rst => false,
    ignore_din_for_gcd => false,
    percent_full_width => 1
  )
  port map (
    en => '1',
    rst => '0',
    din => addsub1_s_net,
    we => constant11_op_net(0),
    re => delay8_q_net(0),
    clk => clk_net,
    ce => ce_net,
    we_ce => ce_net,
    re_ce => ce_net,
    dout => fifo1_dout_net,
    empty => fifo1_empty_net,
    full => fifo1_full_net
  );
  reinterpret1 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => fifo1_dout_net,
    output_port => reinterpret1_output_port_net
  );
end structural;
-- Generated from Simulink block PSB3_0/DPRAM_FIR_Coeffs_1/Scalar to Vector
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_scalar_to_vector is
  port (
    i : in std_logic_vector( 256-1 downto 0 );
    o_1 : out std_logic_vector( 16-1 downto 0 );
    o_2 : out std_logic_vector( 16-1 downto 0 );
    o_3 : out std_logic_vector( 16-1 downto 0 );
    o_4 : out std_logic_vector( 16-1 downto 0 );
    o_5 : out std_logic_vector( 16-1 downto 0 );
    o_6 : out std_logic_vector( 16-1 downto 0 );
    o_7 : out std_logic_vector( 16-1 downto 0 );
    o_8 : out std_logic_vector( 16-1 downto 0 );
    o_9 : out std_logic_vector( 16-1 downto 0 );
    o_10 : out std_logic_vector( 16-1 downto 0 );
    o_11 : out std_logic_vector( 16-1 downto 0 );
    o_12 : out std_logic_vector( 16-1 downto 0 );
    o_13 : out std_logic_vector( 16-1 downto 0 );
    o_14 : out std_logic_vector( 16-1 downto 0 );
    o_15 : out std_logic_vector( 16-1 downto 0 );
    o_16 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_scalar_to_vector;
architecture structural of psb3_0_scalar_to_vector is 
  signal slice1_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 16-1 downto 0 );
  signal dpram_fir_coeffs_1_douta_net : std_logic_vector( 256-1 downto 0 );
begin
  o_1 <= slice0_y_net;
  o_2 <= slice1_y_net;
  o_3 <= slice2_y_net;
  o_4 <= slice3_y_net;
  o_5 <= slice4_y_net;
  o_6 <= slice5_y_net;
  o_7 <= slice6_y_net;
  o_8 <= slice7_y_net;
  o_9 <= slice8_y_net;
  o_10 <= slice9_y_net;
  o_11 <= slice10_y_net;
  o_12 <= slice11_y_net;
  o_13 <= slice12_y_net;
  o_14 <= slice13_y_net;
  o_15 <= slice14_y_net;
  o_16 <= slice15_y_net;
  dpram_fir_coeffs_1_douta_net <= i;
  slice0 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 15,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => dpram_fir_coeffs_1_douta_net,
    y => slice0_y_net
  );
  slice1 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 16,
    new_msb => 31,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => dpram_fir_coeffs_1_douta_net,
    y => slice1_y_net
  );
  slice2 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 32,
    new_msb => 47,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => dpram_fir_coeffs_1_douta_net,
    y => slice2_y_net
  );
  slice3 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 48,
    new_msb => 63,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => dpram_fir_coeffs_1_douta_net,
    y => slice3_y_net
  );
  slice4 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 64,
    new_msb => 79,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => dpram_fir_coeffs_1_douta_net,
    y => slice4_y_net
  );
  slice5 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 80,
    new_msb => 95,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => dpram_fir_coeffs_1_douta_net,
    y => slice5_y_net
  );
  slice6 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 96,
    new_msb => 111,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => dpram_fir_coeffs_1_douta_net,
    y => slice6_y_net
  );
  slice7 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 112,
    new_msb => 127,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => dpram_fir_coeffs_1_douta_net,
    y => slice7_y_net
  );
  slice8 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 128,
    new_msb => 143,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => dpram_fir_coeffs_1_douta_net,
    y => slice8_y_net
  );
  slice9 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 144,
    new_msb => 159,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => dpram_fir_coeffs_1_douta_net,
    y => slice9_y_net
  );
  slice10 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 160,
    new_msb => 175,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => dpram_fir_coeffs_1_douta_net,
    y => slice10_y_net
  );
  slice11 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 176,
    new_msb => 191,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => dpram_fir_coeffs_1_douta_net,
    y => slice11_y_net
  );
  slice12 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 192,
    new_msb => 207,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => dpram_fir_coeffs_1_douta_net,
    y => slice12_y_net
  );
  slice13 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 208,
    new_msb => 223,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => dpram_fir_coeffs_1_douta_net,
    y => slice13_y_net
  );
  slice14 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 224,
    new_msb => 239,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => dpram_fir_coeffs_1_douta_net,
    y => slice14_y_net
  );
  slice15 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 240,
    new_msb => 255,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => dpram_fir_coeffs_1_douta_net,
    y => slice15_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/DPRAM_FIR_Coeffs_1/Vector Reinterpret
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_reinterpret is
  port (
    in_1 : in std_logic_vector( 16-1 downto 0 );
    in_2 : in std_logic_vector( 16-1 downto 0 );
    in_3 : in std_logic_vector( 16-1 downto 0 );
    in_4 : in std_logic_vector( 16-1 downto 0 );
    in_5 : in std_logic_vector( 16-1 downto 0 );
    in_6 : in std_logic_vector( 16-1 downto 0 );
    in_7 : in std_logic_vector( 16-1 downto 0 );
    in_8 : in std_logic_vector( 16-1 downto 0 );
    in_9 : in std_logic_vector( 16-1 downto 0 );
    in_10 : in std_logic_vector( 16-1 downto 0 );
    in_11 : in std_logic_vector( 16-1 downto 0 );
    in_12 : in std_logic_vector( 16-1 downto 0 );
    in_13 : in std_logic_vector( 16-1 downto 0 );
    in_14 : in std_logic_vector( 16-1 downto 0 );
    in_15 : in std_logic_vector( 16-1 downto 0 );
    in_16 : in std_logic_vector( 16-1 downto 0 );
    out_1 : out std_logic_vector( 16-1 downto 0 );
    out_2 : out std_logic_vector( 16-1 downto 0 );
    out_3 : out std_logic_vector( 16-1 downto 0 );
    out_4 : out std_logic_vector( 16-1 downto 0 );
    out_5 : out std_logic_vector( 16-1 downto 0 );
    out_6 : out std_logic_vector( 16-1 downto 0 );
    out_7 : out std_logic_vector( 16-1 downto 0 );
    out_8 : out std_logic_vector( 16-1 downto 0 );
    out_9 : out std_logic_vector( 16-1 downto 0 );
    out_10 : out std_logic_vector( 16-1 downto 0 );
    out_11 : out std_logic_vector( 16-1 downto 0 );
    out_12 : out std_logic_vector( 16-1 downto 0 );
    out_13 : out std_logic_vector( 16-1 downto 0 );
    out_14 : out std_logic_vector( 16-1 downto 0 );
    out_15 : out std_logic_vector( 16-1 downto 0 );
    out_16 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_vector_reinterpret;
architecture structural of psb3_0_vector_reinterpret is 
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 16-1 downto 0 );
begin
  out_1 <= reinterpret0_output_port_net;
  out_2 <= reinterpret1_output_port_net;
  out_3 <= reinterpret2_output_port_net;
  out_4 <= reinterpret3_output_port_net;
  out_5 <= reinterpret4_output_port_net;
  out_6 <= reinterpret5_output_port_net;
  out_7 <= reinterpret6_output_port_net;
  out_8 <= reinterpret7_output_port_net;
  out_9 <= reinterpret8_output_port_net;
  out_10 <= reinterpret9_output_port_net;
  out_11 <= reinterpret10_output_port_net;
  out_12 <= reinterpret11_output_port_net;
  out_13 <= reinterpret12_output_port_net;
  out_14 <= reinterpret13_output_port_net;
  out_15 <= reinterpret14_output_port_net;
  out_16 <= reinterpret15_output_port_net;
  slice0_y_net <= in_1;
  slice1_y_net <= in_2;
  slice2_y_net <= in_3;
  slice3_y_net <= in_4;
  slice4_y_net <= in_5;
  slice5_y_net <= in_6;
  slice6_y_net <= in_7;
  slice7_y_net <= in_8;
  slice8_y_net <= in_9;
  slice9_y_net <= in_10;
  slice10_y_net <= in_11;
  slice11_y_net <= in_12;
  slice12_y_net <= in_13;
  slice13_y_net <= in_14;
  slice14_y_net <= in_15;
  slice15_y_net <= in_16;
  reinterpret0 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice0_y_net,
    output_port => reinterpret0_output_port_net
  );
  reinterpret1 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice1_y_net,
    output_port => reinterpret1_output_port_net
  );
  reinterpret2 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice2_y_net,
    output_port => reinterpret2_output_port_net
  );
  reinterpret3 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice3_y_net,
    output_port => reinterpret3_output_port_net
  );
  reinterpret4 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice4_y_net,
    output_port => reinterpret4_output_port_net
  );
  reinterpret5 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice5_y_net,
    output_port => reinterpret5_output_port_net
  );
  reinterpret6 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice6_y_net,
    output_port => reinterpret6_output_port_net
  );
  reinterpret7 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice7_y_net,
    output_port => reinterpret7_output_port_net
  );
  reinterpret8 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice8_y_net,
    output_port => reinterpret8_output_port_net
  );
  reinterpret9 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice9_y_net,
    output_port => reinterpret9_output_port_net
  );
  reinterpret10 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice10_y_net,
    output_port => reinterpret10_output_port_net
  );
  reinterpret11 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice11_y_net,
    output_port => reinterpret11_output_port_net
  );
  reinterpret12 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice12_y_net,
    output_port => reinterpret12_output_port_net
  );
  reinterpret13 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice13_y_net,
    output_port => reinterpret13_output_port_net
  );
  reinterpret14 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice14_y_net,
    output_port => reinterpret14_output_port_net
  );
  reinterpret15 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice15_y_net,
    output_port => reinterpret15_output_port_net
  );
end structural;
-- Generated from Simulink block PSB3_0/DPRAM_FIR_Coeffs_1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_dpram_fir_coeffs_1 is
  port (
    in_rst : in std_logic_vector( 1-1 downto 0 );
    in_en : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    out_fir_coeffs_1 : out std_logic_vector( 16-1 downto 0 );
    out_fir_coeffs_2 : out std_logic_vector( 16-1 downto 0 );
    out_fir_coeffs_3 : out std_logic_vector( 16-1 downto 0 );
    out_fir_coeffs_4 : out std_logic_vector( 16-1 downto 0 );
    out_fir_coeffs_5 : out std_logic_vector( 16-1 downto 0 );
    out_fir_coeffs_6 : out std_logic_vector( 16-1 downto 0 );
    out_fir_coeffs_7 : out std_logic_vector( 16-1 downto 0 );
    out_fir_coeffs_8 : out std_logic_vector( 16-1 downto 0 );
    out_fir_coeffs_9 : out std_logic_vector( 16-1 downto 0 );
    out_fir_coeffs_10 : out std_logic_vector( 16-1 downto 0 );
    out_fir_coeffs_11 : out std_logic_vector( 16-1 downto 0 );
    out_fir_coeffs_12 : out std_logic_vector( 16-1 downto 0 );
    out_fir_coeffs_13 : out std_logic_vector( 16-1 downto 0 );
    out_fir_coeffs_14 : out std_logic_vector( 16-1 downto 0 );
    out_fir_coeffs_15 : out std_logic_vector( 16-1 downto 0 );
    out_fir_coeffs_16 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_dpram_fir_coeffs_1;
architecture structural of psb3_0_dpram_fir_coeffs_1 is 
  signal dpram_fir_coeffs_1_doutb_net : std_logic_vector( 256-1 downto 0 );
  signal read_addr_op_net : std_logic_vector( 8-1 downto 0 );
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal clk_net : std_logic;
  signal ce_net : std_logic;
  signal slice0_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 16-1 downto 0 );
  signal gin_tl_reset_net : std_logic_vector( 1-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 16-1 downto 0 );
  signal constant2_op_net : std_logic_vector( 1-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 16-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 256-1 downto 0 );
  signal dpram_fir_coeffs_1_douta_net : std_logic_vector( 256-1 downto 0 );
  signal constant0_op_net : std_logic_vector( 8-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 16-1 downto 0 );
begin
  out_fir_coeffs_1 <= reinterpret0_output_port_net;
  out_fir_coeffs_2 <= reinterpret1_output_port_net;
  out_fir_coeffs_3 <= reinterpret2_output_port_net;
  out_fir_coeffs_4 <= reinterpret3_output_port_net;
  out_fir_coeffs_5 <= reinterpret4_output_port_net;
  out_fir_coeffs_6 <= reinterpret5_output_port_net;
  out_fir_coeffs_7 <= reinterpret6_output_port_net;
  out_fir_coeffs_8 <= reinterpret7_output_port_net;
  out_fir_coeffs_9 <= reinterpret8_output_port_net;
  out_fir_coeffs_10 <= reinterpret9_output_port_net;
  out_fir_coeffs_11 <= reinterpret10_output_port_net;
  out_fir_coeffs_12 <= reinterpret11_output_port_net;
  out_fir_coeffs_13 <= reinterpret12_output_port_net;
  out_fir_coeffs_14 <= reinterpret13_output_port_net;
  out_fir_coeffs_15 <= reinterpret14_output_port_net;
  out_fir_coeffs_16 <= reinterpret15_output_port_net;
  gin_tl_reset_net <= in_rst;
  delay8_q_net <= in_en;
  clk_net <= clk_1;
  ce_net <= ce_1;
  scalar_to_vector : entity xil_defaultlib.psb3_0_scalar_to_vector 
  port map (
    i => dpram_fir_coeffs_1_douta_net,
    o_1 => slice0_y_net,
    o_2 => slice1_y_net,
    o_3 => slice2_y_net,
    o_4 => slice3_y_net,
    o_5 => slice4_y_net,
    o_6 => slice5_y_net,
    o_7 => slice6_y_net,
    o_8 => slice7_y_net,
    o_9 => slice8_y_net,
    o_10 => slice9_y_net,
    o_11 => slice10_y_net,
    o_12 => slice11_y_net,
    o_13 => slice12_y_net,
    o_14 => slice13_y_net,
    o_15 => slice14_y_net,
    o_16 => slice15_y_net
  );
  vector_reinterpret : entity xil_defaultlib.psb3_0_vector_reinterpret 
  port map (
    in_1 => slice0_y_net,
    in_2 => slice1_y_net,
    in_3 => slice2_y_net,
    in_4 => slice3_y_net,
    in_5 => slice4_y_net,
    in_6 => slice5_y_net,
    in_7 => slice6_y_net,
    in_8 => slice7_y_net,
    in_9 => slice8_y_net,
    in_10 => slice9_y_net,
    in_11 => slice10_y_net,
    in_12 => slice11_y_net,
    in_13 => slice12_y_net,
    in_14 => slice13_y_net,
    in_15 => slice14_y_net,
    in_16 => slice15_y_net,
    out_1 => reinterpret0_output_port_net,
    out_2 => reinterpret1_output_port_net,
    out_3 => reinterpret2_output_port_net,
    out_4 => reinterpret3_output_port_net,
    out_5 => reinterpret4_output_port_net,
    out_6 => reinterpret5_output_port_net,
    out_7 => reinterpret6_output_port_net,
    out_8 => reinterpret7_output_port_net,
    out_9 => reinterpret8_output_port_net,
    out_10 => reinterpret9_output_port_net,
    out_11 => reinterpret10_output_port_net,
    out_12 => reinterpret11_output_port_net,
    out_13 => reinterpret12_output_port_net,
    out_14 => reinterpret13_output_port_net,
    out_15 => reinterpret14_output_port_net,
    out_16 => reinterpret15_output_port_net
  );
  constant0 : entity xil_defaultlib.sysgen_constant_0714509e7f 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant0_op_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_31aefdfd97 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  constant2 : entity xil_defaultlib.sysgen_constant_de9059c03f 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant2_op_net
  );
  dpram_fir_coeffs_1 : entity xil_defaultlib.psb3_0_xltdpram 
  generic map (
    addr_width_b => 8,
    clocking_mode => "common_clock",
    data_width_b => 256,
    latency => 2,
    mem_init_file => "xpm_6cc9b6_vivado.mem",
    mem_size => 65536,
    mem_type => "block",
    read_reset_a => "0",
    read_reset_b => "0",
    width => 256,
    width_addr => 8,
    write_mode_a => "no_change",
    write_mode_b => "no_change"
  )
  port map (
    ena => "1",
    enb => "1",
    rsta => "0",
    rstb => "0",
    addra => read_addr_op_net,
    dina => constant1_op_net,
    wea => constant2_op_net,
    addrb => constant0_op_net,
    dinb => constant1_op_net,
    web => constant2_op_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dpram_fir_coeffs_1_douta_net,
    doutb => dpram_fir_coeffs_1_doutb_net
  );
  read_addr : entity xil_defaultlib.psb3_0_xlcounter_free 
  generic map (
    core_name0 => "psb3_0_c_counter_binary_v12_0_i0",
    op_arith => xlUnsigned,
    op_width => 8
  )
  port map (
    clr => '0',
    rst => gin_tl_reset_net,
    en => delay8_q_net,
    clk => clk_net,
    ce => ce_net,
    op => read_addr_op_net
  );
end structural;
-- Generated from Simulink block PSB3_0/DPRAM_FIR_Coeffs_2/Scalar to Vector
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_scalar_to_vector_x0 is
  port (
    i : in std_logic_vector( 256-1 downto 0 );
    o_1 : out std_logic_vector( 16-1 downto 0 );
    o_2 : out std_logic_vector( 16-1 downto 0 );
    o_3 : out std_logic_vector( 16-1 downto 0 );
    o_4 : out std_logic_vector( 16-1 downto 0 );
    o_5 : out std_logic_vector( 16-1 downto 0 );
    o_6 : out std_logic_vector( 16-1 downto 0 );
    o_7 : out std_logic_vector( 16-1 downto 0 );
    o_8 : out std_logic_vector( 16-1 downto 0 );
    o_9 : out std_logic_vector( 16-1 downto 0 );
    o_10 : out std_logic_vector( 16-1 downto 0 );
    o_11 : out std_logic_vector( 16-1 downto 0 );
    o_12 : out std_logic_vector( 16-1 downto 0 );
    o_13 : out std_logic_vector( 16-1 downto 0 );
    o_14 : out std_logic_vector( 16-1 downto 0 );
    o_15 : out std_logic_vector( 16-1 downto 0 );
    o_16 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_scalar_to_vector_x0;
architecture structural of psb3_0_scalar_to_vector_x0 is 
  signal slice15_y_net : std_logic_vector( 16-1 downto 0 );
  signal dpram_fir_coeffs_2_douta_net : std_logic_vector( 256-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 16-1 downto 0 );
begin
  o_1 <= slice0_y_net;
  o_2 <= slice1_y_net;
  o_3 <= slice2_y_net;
  o_4 <= slice3_y_net;
  o_5 <= slice4_y_net;
  o_6 <= slice5_y_net;
  o_7 <= slice6_y_net;
  o_8 <= slice7_y_net;
  o_9 <= slice8_y_net;
  o_10 <= slice9_y_net;
  o_11 <= slice10_y_net;
  o_12 <= slice11_y_net;
  o_13 <= slice12_y_net;
  o_14 <= slice13_y_net;
  o_15 <= slice14_y_net;
  o_16 <= slice15_y_net;
  dpram_fir_coeffs_2_douta_net <= i;
  slice0 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 15,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => dpram_fir_coeffs_2_douta_net,
    y => slice0_y_net
  );
  slice1 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 16,
    new_msb => 31,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => dpram_fir_coeffs_2_douta_net,
    y => slice1_y_net
  );
  slice2 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 32,
    new_msb => 47,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => dpram_fir_coeffs_2_douta_net,
    y => slice2_y_net
  );
  slice3 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 48,
    new_msb => 63,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => dpram_fir_coeffs_2_douta_net,
    y => slice3_y_net
  );
  slice4 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 64,
    new_msb => 79,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => dpram_fir_coeffs_2_douta_net,
    y => slice4_y_net
  );
  slice5 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 80,
    new_msb => 95,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => dpram_fir_coeffs_2_douta_net,
    y => slice5_y_net
  );
  slice6 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 96,
    new_msb => 111,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => dpram_fir_coeffs_2_douta_net,
    y => slice6_y_net
  );
  slice7 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 112,
    new_msb => 127,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => dpram_fir_coeffs_2_douta_net,
    y => slice7_y_net
  );
  slice8 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 128,
    new_msb => 143,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => dpram_fir_coeffs_2_douta_net,
    y => slice8_y_net
  );
  slice9 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 144,
    new_msb => 159,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => dpram_fir_coeffs_2_douta_net,
    y => slice9_y_net
  );
  slice10 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 160,
    new_msb => 175,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => dpram_fir_coeffs_2_douta_net,
    y => slice10_y_net
  );
  slice11 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 176,
    new_msb => 191,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => dpram_fir_coeffs_2_douta_net,
    y => slice11_y_net
  );
  slice12 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 192,
    new_msb => 207,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => dpram_fir_coeffs_2_douta_net,
    y => slice12_y_net
  );
  slice13 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 208,
    new_msb => 223,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => dpram_fir_coeffs_2_douta_net,
    y => slice13_y_net
  );
  slice14 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 224,
    new_msb => 239,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => dpram_fir_coeffs_2_douta_net,
    y => slice14_y_net
  );
  slice15 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 240,
    new_msb => 255,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => dpram_fir_coeffs_2_douta_net,
    y => slice15_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/DPRAM_FIR_Coeffs_2/Vector Reinterpret
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_reinterpret_x0 is
  port (
    in_1 : in std_logic_vector( 16-1 downto 0 );
    in_2 : in std_logic_vector( 16-1 downto 0 );
    in_3 : in std_logic_vector( 16-1 downto 0 );
    in_4 : in std_logic_vector( 16-1 downto 0 );
    in_5 : in std_logic_vector( 16-1 downto 0 );
    in_6 : in std_logic_vector( 16-1 downto 0 );
    in_7 : in std_logic_vector( 16-1 downto 0 );
    in_8 : in std_logic_vector( 16-1 downto 0 );
    in_9 : in std_logic_vector( 16-1 downto 0 );
    in_10 : in std_logic_vector( 16-1 downto 0 );
    in_11 : in std_logic_vector( 16-1 downto 0 );
    in_12 : in std_logic_vector( 16-1 downto 0 );
    in_13 : in std_logic_vector( 16-1 downto 0 );
    in_14 : in std_logic_vector( 16-1 downto 0 );
    in_15 : in std_logic_vector( 16-1 downto 0 );
    in_16 : in std_logic_vector( 16-1 downto 0 );
    out_1 : out std_logic_vector( 16-1 downto 0 );
    out_2 : out std_logic_vector( 16-1 downto 0 );
    out_3 : out std_logic_vector( 16-1 downto 0 );
    out_4 : out std_logic_vector( 16-1 downto 0 );
    out_5 : out std_logic_vector( 16-1 downto 0 );
    out_6 : out std_logic_vector( 16-1 downto 0 );
    out_7 : out std_logic_vector( 16-1 downto 0 );
    out_8 : out std_logic_vector( 16-1 downto 0 );
    out_9 : out std_logic_vector( 16-1 downto 0 );
    out_10 : out std_logic_vector( 16-1 downto 0 );
    out_11 : out std_logic_vector( 16-1 downto 0 );
    out_12 : out std_logic_vector( 16-1 downto 0 );
    out_13 : out std_logic_vector( 16-1 downto 0 );
    out_14 : out std_logic_vector( 16-1 downto 0 );
    out_15 : out std_logic_vector( 16-1 downto 0 );
    out_16 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_vector_reinterpret_x0;
architecture structural of psb3_0_vector_reinterpret_x0 is 
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 16-1 downto 0 );
begin
  out_1 <= reinterpret0_output_port_net;
  out_2 <= reinterpret1_output_port_net;
  out_3 <= reinterpret2_output_port_net;
  out_4 <= reinterpret3_output_port_net;
  out_5 <= reinterpret4_output_port_net;
  out_6 <= reinterpret5_output_port_net;
  out_7 <= reinterpret6_output_port_net;
  out_8 <= reinterpret7_output_port_net;
  out_9 <= reinterpret8_output_port_net;
  out_10 <= reinterpret9_output_port_net;
  out_11 <= reinterpret10_output_port_net;
  out_12 <= reinterpret11_output_port_net;
  out_13 <= reinterpret12_output_port_net;
  out_14 <= reinterpret13_output_port_net;
  out_15 <= reinterpret14_output_port_net;
  out_16 <= reinterpret15_output_port_net;
  slice0_y_net <= in_1;
  slice1_y_net <= in_2;
  slice2_y_net <= in_3;
  slice3_y_net <= in_4;
  slice4_y_net <= in_5;
  slice5_y_net <= in_6;
  slice6_y_net <= in_7;
  slice7_y_net <= in_8;
  slice8_y_net <= in_9;
  slice9_y_net <= in_10;
  slice10_y_net <= in_11;
  slice11_y_net <= in_12;
  slice12_y_net <= in_13;
  slice13_y_net <= in_14;
  slice14_y_net <= in_15;
  slice15_y_net <= in_16;
  reinterpret0 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice0_y_net,
    output_port => reinterpret0_output_port_net
  );
  reinterpret1 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice1_y_net,
    output_port => reinterpret1_output_port_net
  );
  reinterpret2 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice2_y_net,
    output_port => reinterpret2_output_port_net
  );
  reinterpret3 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice3_y_net,
    output_port => reinterpret3_output_port_net
  );
  reinterpret4 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice4_y_net,
    output_port => reinterpret4_output_port_net
  );
  reinterpret5 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice5_y_net,
    output_port => reinterpret5_output_port_net
  );
  reinterpret6 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice6_y_net,
    output_port => reinterpret6_output_port_net
  );
  reinterpret7 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice7_y_net,
    output_port => reinterpret7_output_port_net
  );
  reinterpret8 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice8_y_net,
    output_port => reinterpret8_output_port_net
  );
  reinterpret9 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice9_y_net,
    output_port => reinterpret9_output_port_net
  );
  reinterpret10 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice10_y_net,
    output_port => reinterpret10_output_port_net
  );
  reinterpret11 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice11_y_net,
    output_port => reinterpret11_output_port_net
  );
  reinterpret12 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice12_y_net,
    output_port => reinterpret12_output_port_net
  );
  reinterpret13 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice13_y_net,
    output_port => reinterpret13_output_port_net
  );
  reinterpret14 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice14_y_net,
    output_port => reinterpret14_output_port_net
  );
  reinterpret15 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice15_y_net,
    output_port => reinterpret15_output_port_net
  );
end structural;
-- Generated from Simulink block PSB3_0/DPRAM_FIR_Coeffs_2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_dpram_fir_coeffs_2 is
  port (
    in_rst : in std_logic_vector( 1-1 downto 0 );
    in_en : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    out_fir_coeffs_1 : out std_logic_vector( 16-1 downto 0 );
    out_fir_coeffs_2 : out std_logic_vector( 16-1 downto 0 );
    out_fir_coeffs_3 : out std_logic_vector( 16-1 downto 0 );
    out_fir_coeffs_4 : out std_logic_vector( 16-1 downto 0 );
    out_fir_coeffs_5 : out std_logic_vector( 16-1 downto 0 );
    out_fir_coeffs_6 : out std_logic_vector( 16-1 downto 0 );
    out_fir_coeffs_7 : out std_logic_vector( 16-1 downto 0 );
    out_fir_coeffs_8 : out std_logic_vector( 16-1 downto 0 );
    out_fir_coeffs_9 : out std_logic_vector( 16-1 downto 0 );
    out_fir_coeffs_10 : out std_logic_vector( 16-1 downto 0 );
    out_fir_coeffs_11 : out std_logic_vector( 16-1 downto 0 );
    out_fir_coeffs_12 : out std_logic_vector( 16-1 downto 0 );
    out_fir_coeffs_13 : out std_logic_vector( 16-1 downto 0 );
    out_fir_coeffs_14 : out std_logic_vector( 16-1 downto 0 );
    out_fir_coeffs_15 : out std_logic_vector( 16-1 downto 0 );
    out_fir_coeffs_16 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_dpram_fir_coeffs_2;
architecture structural of psb3_0_dpram_fir_coeffs_2 is 
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal gin_tl_reset_net : std_logic_vector( 1-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 16-1 downto 0 );
  signal ce_net : std_logic;
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal clk_net : std_logic;
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 16-1 downto 0 );
  signal dpram_fir_coeffs_2_douta_net : std_logic_vector( 256-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal constant2_op_net : std_logic_vector( 1-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 256-1 downto 0 );
  signal read_addr_op_net : std_logic_vector( 8-1 downto 0 );
  signal dpram_fir_coeffs_2_doutb_net : std_logic_vector( 256-1 downto 0 );
  signal constant0_op_net : std_logic_vector( 8-1 downto 0 );
begin
  out_fir_coeffs_1 <= reinterpret0_output_port_net;
  out_fir_coeffs_2 <= reinterpret1_output_port_net;
  out_fir_coeffs_3 <= reinterpret2_output_port_net;
  out_fir_coeffs_4 <= reinterpret3_output_port_net;
  out_fir_coeffs_5 <= reinterpret4_output_port_net;
  out_fir_coeffs_6 <= reinterpret5_output_port_net;
  out_fir_coeffs_7 <= reinterpret6_output_port_net;
  out_fir_coeffs_8 <= reinterpret7_output_port_net;
  out_fir_coeffs_9 <= reinterpret8_output_port_net;
  out_fir_coeffs_10 <= reinterpret9_output_port_net;
  out_fir_coeffs_11 <= reinterpret10_output_port_net;
  out_fir_coeffs_12 <= reinterpret11_output_port_net;
  out_fir_coeffs_13 <= reinterpret12_output_port_net;
  out_fir_coeffs_14 <= reinterpret13_output_port_net;
  out_fir_coeffs_15 <= reinterpret14_output_port_net;
  out_fir_coeffs_16 <= reinterpret15_output_port_net;
  gin_tl_reset_net <= in_rst;
  delay8_q_net <= in_en;
  clk_net <= clk_1;
  ce_net <= ce_1;
  scalar_to_vector : entity xil_defaultlib.psb3_0_scalar_to_vector_x0 
  port map (
    i => dpram_fir_coeffs_2_douta_net,
    o_1 => slice0_y_net,
    o_2 => slice1_y_net,
    o_3 => slice2_y_net,
    o_4 => slice3_y_net,
    o_5 => slice4_y_net,
    o_6 => slice5_y_net,
    o_7 => slice6_y_net,
    o_8 => slice7_y_net,
    o_9 => slice8_y_net,
    o_10 => slice9_y_net,
    o_11 => slice10_y_net,
    o_12 => slice11_y_net,
    o_13 => slice12_y_net,
    o_14 => slice13_y_net,
    o_15 => slice14_y_net,
    o_16 => slice15_y_net
  );
  vector_reinterpret : entity xil_defaultlib.psb3_0_vector_reinterpret_x0 
  port map (
    in_1 => slice0_y_net,
    in_2 => slice1_y_net,
    in_3 => slice2_y_net,
    in_4 => slice3_y_net,
    in_5 => slice4_y_net,
    in_6 => slice5_y_net,
    in_7 => slice6_y_net,
    in_8 => slice7_y_net,
    in_9 => slice8_y_net,
    in_10 => slice9_y_net,
    in_11 => slice10_y_net,
    in_12 => slice11_y_net,
    in_13 => slice12_y_net,
    in_14 => slice13_y_net,
    in_15 => slice14_y_net,
    in_16 => slice15_y_net,
    out_1 => reinterpret0_output_port_net,
    out_2 => reinterpret1_output_port_net,
    out_3 => reinterpret2_output_port_net,
    out_4 => reinterpret3_output_port_net,
    out_5 => reinterpret4_output_port_net,
    out_6 => reinterpret5_output_port_net,
    out_7 => reinterpret6_output_port_net,
    out_8 => reinterpret7_output_port_net,
    out_9 => reinterpret8_output_port_net,
    out_10 => reinterpret9_output_port_net,
    out_11 => reinterpret10_output_port_net,
    out_12 => reinterpret11_output_port_net,
    out_13 => reinterpret12_output_port_net,
    out_14 => reinterpret13_output_port_net,
    out_15 => reinterpret14_output_port_net,
    out_16 => reinterpret15_output_port_net
  );
  constant0 : entity xil_defaultlib.sysgen_constant_0714509e7f 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant0_op_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_31aefdfd97 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  constant2 : entity xil_defaultlib.sysgen_constant_de9059c03f 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant2_op_net
  );
  dpram_fir_coeffs_2 : entity xil_defaultlib.psb3_0_xltdpram 
  generic map (
    addr_width_b => 8,
    clocking_mode => "common_clock",
    data_width_b => 256,
    latency => 2,
    mem_init_file => "xpm_5d2d2a_vivado.mem",
    mem_size => 65536,
    mem_type => "block",
    read_reset_a => "0",
    read_reset_b => "0",
    width => 256,
    width_addr => 8,
    write_mode_a => "no_change",
    write_mode_b => "no_change"
  )
  port map (
    ena => "1",
    enb => "1",
    rsta => "0",
    rstb => "0",
    addra => read_addr_op_net,
    dina => constant1_op_net,
    wea => constant2_op_net,
    addrb => constant0_op_net,
    dinb => constant1_op_net,
    web => constant2_op_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dpram_fir_coeffs_2_douta_net,
    doutb => dpram_fir_coeffs_2_doutb_net
  );
  read_addr : entity xil_defaultlib.psb3_0_xlcounter_free 
  generic map (
    core_name0 => "psb3_0_c_counter_binary_v12_0_i0",
    op_arith => xlUnsigned,
    op_width => 8
  )
  port map (
    clr => '0',
    rst => gin_tl_reset_net,
    en => delay8_q_net,
    clk => clk_net,
    ce => ce_net,
    op => read_addr_op_net
  );
end structural;
-- Generated from Simulink block PSB3_0/DPRAM_FIR_Coeffs_3/Scalar to Vector
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_scalar_to_vector_x1 is
  port (
    i : in std_logic_vector( 256-1 downto 0 );
    o_1 : out std_logic_vector( 16-1 downto 0 );
    o_2 : out std_logic_vector( 16-1 downto 0 );
    o_3 : out std_logic_vector( 16-1 downto 0 );
    o_4 : out std_logic_vector( 16-1 downto 0 );
    o_5 : out std_logic_vector( 16-1 downto 0 );
    o_6 : out std_logic_vector( 16-1 downto 0 );
    o_7 : out std_logic_vector( 16-1 downto 0 );
    o_8 : out std_logic_vector( 16-1 downto 0 );
    o_9 : out std_logic_vector( 16-1 downto 0 );
    o_10 : out std_logic_vector( 16-1 downto 0 );
    o_11 : out std_logic_vector( 16-1 downto 0 );
    o_12 : out std_logic_vector( 16-1 downto 0 );
    o_13 : out std_logic_vector( 16-1 downto 0 );
    o_14 : out std_logic_vector( 16-1 downto 0 );
    o_15 : out std_logic_vector( 16-1 downto 0 );
    o_16 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_scalar_to_vector_x1;
architecture structural of psb3_0_scalar_to_vector_x1 is 
  signal slice1_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 16-1 downto 0 );
  signal dpram_fir_coeffs_3_douta_net : std_logic_vector( 256-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 16-1 downto 0 );
begin
  o_1 <= slice0_y_net;
  o_2 <= slice1_y_net;
  o_3 <= slice2_y_net;
  o_4 <= slice3_y_net;
  o_5 <= slice4_y_net;
  o_6 <= slice5_y_net;
  o_7 <= slice6_y_net;
  o_8 <= slice7_y_net;
  o_9 <= slice8_y_net;
  o_10 <= slice9_y_net;
  o_11 <= slice10_y_net;
  o_12 <= slice11_y_net;
  o_13 <= slice12_y_net;
  o_14 <= slice13_y_net;
  o_15 <= slice14_y_net;
  o_16 <= slice15_y_net;
  dpram_fir_coeffs_3_douta_net <= i;
  slice0 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 15,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => dpram_fir_coeffs_3_douta_net,
    y => slice0_y_net
  );
  slice1 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 16,
    new_msb => 31,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => dpram_fir_coeffs_3_douta_net,
    y => slice1_y_net
  );
  slice2 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 32,
    new_msb => 47,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => dpram_fir_coeffs_3_douta_net,
    y => slice2_y_net
  );
  slice3 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 48,
    new_msb => 63,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => dpram_fir_coeffs_3_douta_net,
    y => slice3_y_net
  );
  slice4 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 64,
    new_msb => 79,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => dpram_fir_coeffs_3_douta_net,
    y => slice4_y_net
  );
  slice5 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 80,
    new_msb => 95,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => dpram_fir_coeffs_3_douta_net,
    y => slice5_y_net
  );
  slice6 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 96,
    new_msb => 111,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => dpram_fir_coeffs_3_douta_net,
    y => slice6_y_net
  );
  slice7 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 112,
    new_msb => 127,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => dpram_fir_coeffs_3_douta_net,
    y => slice7_y_net
  );
  slice8 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 128,
    new_msb => 143,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => dpram_fir_coeffs_3_douta_net,
    y => slice8_y_net
  );
  slice9 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 144,
    new_msb => 159,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => dpram_fir_coeffs_3_douta_net,
    y => slice9_y_net
  );
  slice10 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 160,
    new_msb => 175,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => dpram_fir_coeffs_3_douta_net,
    y => slice10_y_net
  );
  slice11 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 176,
    new_msb => 191,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => dpram_fir_coeffs_3_douta_net,
    y => slice11_y_net
  );
  slice12 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 192,
    new_msb => 207,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => dpram_fir_coeffs_3_douta_net,
    y => slice12_y_net
  );
  slice13 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 208,
    new_msb => 223,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => dpram_fir_coeffs_3_douta_net,
    y => slice13_y_net
  );
  slice14 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 224,
    new_msb => 239,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => dpram_fir_coeffs_3_douta_net,
    y => slice14_y_net
  );
  slice15 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 240,
    new_msb => 255,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => dpram_fir_coeffs_3_douta_net,
    y => slice15_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/DPRAM_FIR_Coeffs_3/Vector Reinterpret
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_reinterpret_x1 is
  port (
    in_1 : in std_logic_vector( 16-1 downto 0 );
    in_2 : in std_logic_vector( 16-1 downto 0 );
    in_3 : in std_logic_vector( 16-1 downto 0 );
    in_4 : in std_logic_vector( 16-1 downto 0 );
    in_5 : in std_logic_vector( 16-1 downto 0 );
    in_6 : in std_logic_vector( 16-1 downto 0 );
    in_7 : in std_logic_vector( 16-1 downto 0 );
    in_8 : in std_logic_vector( 16-1 downto 0 );
    in_9 : in std_logic_vector( 16-1 downto 0 );
    in_10 : in std_logic_vector( 16-1 downto 0 );
    in_11 : in std_logic_vector( 16-1 downto 0 );
    in_12 : in std_logic_vector( 16-1 downto 0 );
    in_13 : in std_logic_vector( 16-1 downto 0 );
    in_14 : in std_logic_vector( 16-1 downto 0 );
    in_15 : in std_logic_vector( 16-1 downto 0 );
    in_16 : in std_logic_vector( 16-1 downto 0 );
    out_1 : out std_logic_vector( 16-1 downto 0 );
    out_2 : out std_logic_vector( 16-1 downto 0 );
    out_3 : out std_logic_vector( 16-1 downto 0 );
    out_4 : out std_logic_vector( 16-1 downto 0 );
    out_5 : out std_logic_vector( 16-1 downto 0 );
    out_6 : out std_logic_vector( 16-1 downto 0 );
    out_7 : out std_logic_vector( 16-1 downto 0 );
    out_8 : out std_logic_vector( 16-1 downto 0 );
    out_9 : out std_logic_vector( 16-1 downto 0 );
    out_10 : out std_logic_vector( 16-1 downto 0 );
    out_11 : out std_logic_vector( 16-1 downto 0 );
    out_12 : out std_logic_vector( 16-1 downto 0 );
    out_13 : out std_logic_vector( 16-1 downto 0 );
    out_14 : out std_logic_vector( 16-1 downto 0 );
    out_15 : out std_logic_vector( 16-1 downto 0 );
    out_16 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_vector_reinterpret_x1;
architecture structural of psb3_0_vector_reinterpret_x1 is 
  signal slice15_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
begin
  out_1 <= reinterpret0_output_port_net;
  out_2 <= reinterpret1_output_port_net;
  out_3 <= reinterpret2_output_port_net;
  out_4 <= reinterpret3_output_port_net;
  out_5 <= reinterpret4_output_port_net;
  out_6 <= reinterpret5_output_port_net;
  out_7 <= reinterpret6_output_port_net;
  out_8 <= reinterpret7_output_port_net;
  out_9 <= reinterpret8_output_port_net;
  out_10 <= reinterpret9_output_port_net;
  out_11 <= reinterpret10_output_port_net;
  out_12 <= reinterpret11_output_port_net;
  out_13 <= reinterpret12_output_port_net;
  out_14 <= reinterpret13_output_port_net;
  out_15 <= reinterpret14_output_port_net;
  out_16 <= reinterpret15_output_port_net;
  slice0_y_net <= in_1;
  slice1_y_net <= in_2;
  slice2_y_net <= in_3;
  slice3_y_net <= in_4;
  slice4_y_net <= in_5;
  slice5_y_net <= in_6;
  slice6_y_net <= in_7;
  slice7_y_net <= in_8;
  slice8_y_net <= in_9;
  slice9_y_net <= in_10;
  slice10_y_net <= in_11;
  slice11_y_net <= in_12;
  slice12_y_net <= in_13;
  slice13_y_net <= in_14;
  slice14_y_net <= in_15;
  slice15_y_net <= in_16;
  reinterpret0 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice0_y_net,
    output_port => reinterpret0_output_port_net
  );
  reinterpret1 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice1_y_net,
    output_port => reinterpret1_output_port_net
  );
  reinterpret2 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice2_y_net,
    output_port => reinterpret2_output_port_net
  );
  reinterpret3 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice3_y_net,
    output_port => reinterpret3_output_port_net
  );
  reinterpret4 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice4_y_net,
    output_port => reinterpret4_output_port_net
  );
  reinterpret5 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice5_y_net,
    output_port => reinterpret5_output_port_net
  );
  reinterpret6 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice6_y_net,
    output_port => reinterpret6_output_port_net
  );
  reinterpret7 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice7_y_net,
    output_port => reinterpret7_output_port_net
  );
  reinterpret8 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice8_y_net,
    output_port => reinterpret8_output_port_net
  );
  reinterpret9 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice9_y_net,
    output_port => reinterpret9_output_port_net
  );
  reinterpret10 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice10_y_net,
    output_port => reinterpret10_output_port_net
  );
  reinterpret11 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice11_y_net,
    output_port => reinterpret11_output_port_net
  );
  reinterpret12 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice12_y_net,
    output_port => reinterpret12_output_port_net
  );
  reinterpret13 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice13_y_net,
    output_port => reinterpret13_output_port_net
  );
  reinterpret14 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice14_y_net,
    output_port => reinterpret14_output_port_net
  );
  reinterpret15 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice15_y_net,
    output_port => reinterpret15_output_port_net
  );
end structural;
-- Generated from Simulink block PSB3_0/DPRAM_FIR_Coeffs_3
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_dpram_fir_coeffs_3 is
  port (
    in_rst : in std_logic_vector( 1-1 downto 0 );
    in_en : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    out_fir_coeffs_1 : out std_logic_vector( 16-1 downto 0 );
    out_fir_coeffs_2 : out std_logic_vector( 16-1 downto 0 );
    out_fir_coeffs_3 : out std_logic_vector( 16-1 downto 0 );
    out_fir_coeffs_4 : out std_logic_vector( 16-1 downto 0 );
    out_fir_coeffs_5 : out std_logic_vector( 16-1 downto 0 );
    out_fir_coeffs_6 : out std_logic_vector( 16-1 downto 0 );
    out_fir_coeffs_7 : out std_logic_vector( 16-1 downto 0 );
    out_fir_coeffs_8 : out std_logic_vector( 16-1 downto 0 );
    out_fir_coeffs_9 : out std_logic_vector( 16-1 downto 0 );
    out_fir_coeffs_10 : out std_logic_vector( 16-1 downto 0 );
    out_fir_coeffs_11 : out std_logic_vector( 16-1 downto 0 );
    out_fir_coeffs_12 : out std_logic_vector( 16-1 downto 0 );
    out_fir_coeffs_13 : out std_logic_vector( 16-1 downto 0 );
    out_fir_coeffs_14 : out std_logic_vector( 16-1 downto 0 );
    out_fir_coeffs_15 : out std_logic_vector( 16-1 downto 0 );
    out_fir_coeffs_16 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_dpram_fir_coeffs_3;
architecture structural of psb3_0_dpram_fir_coeffs_3 is 
  signal dpram_fir_coeffs_3_doutb_net : std_logic_vector( 256-1 downto 0 );
  signal read_addr_op_net : std_logic_vector( 8-1 downto 0 );
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal clk_net : std_logic;
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal ce_net : std_logic;
  signal slice1_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal gin_tl_reset_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal constant2_op_net : std_logic_vector( 1-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 16-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 256-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 16-1 downto 0 );
  signal constant0_op_net : std_logic_vector( 8-1 downto 0 );
  signal dpram_fir_coeffs_3_douta_net : std_logic_vector( 256-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 16-1 downto 0 );
begin
  out_fir_coeffs_1 <= reinterpret0_output_port_net;
  out_fir_coeffs_2 <= reinterpret1_output_port_net;
  out_fir_coeffs_3 <= reinterpret2_output_port_net;
  out_fir_coeffs_4 <= reinterpret3_output_port_net;
  out_fir_coeffs_5 <= reinterpret4_output_port_net;
  out_fir_coeffs_6 <= reinterpret5_output_port_net;
  out_fir_coeffs_7 <= reinterpret6_output_port_net;
  out_fir_coeffs_8 <= reinterpret7_output_port_net;
  out_fir_coeffs_9 <= reinterpret8_output_port_net;
  out_fir_coeffs_10 <= reinterpret9_output_port_net;
  out_fir_coeffs_11 <= reinterpret10_output_port_net;
  out_fir_coeffs_12 <= reinterpret11_output_port_net;
  out_fir_coeffs_13 <= reinterpret12_output_port_net;
  out_fir_coeffs_14 <= reinterpret13_output_port_net;
  out_fir_coeffs_15 <= reinterpret14_output_port_net;
  out_fir_coeffs_16 <= reinterpret15_output_port_net;
  gin_tl_reset_net <= in_rst;
  delay8_q_net <= in_en;
  clk_net <= clk_1;
  ce_net <= ce_1;
  scalar_to_vector : entity xil_defaultlib.psb3_0_scalar_to_vector_x1 
  port map (
    i => dpram_fir_coeffs_3_douta_net,
    o_1 => slice0_y_net,
    o_2 => slice1_y_net,
    o_3 => slice2_y_net,
    o_4 => slice3_y_net,
    o_5 => slice4_y_net,
    o_6 => slice5_y_net,
    o_7 => slice6_y_net,
    o_8 => slice7_y_net,
    o_9 => slice8_y_net,
    o_10 => slice9_y_net,
    o_11 => slice10_y_net,
    o_12 => slice11_y_net,
    o_13 => slice12_y_net,
    o_14 => slice13_y_net,
    o_15 => slice14_y_net,
    o_16 => slice15_y_net
  );
  vector_reinterpret : entity xil_defaultlib.psb3_0_vector_reinterpret_x1 
  port map (
    in_1 => slice0_y_net,
    in_2 => slice1_y_net,
    in_3 => slice2_y_net,
    in_4 => slice3_y_net,
    in_5 => slice4_y_net,
    in_6 => slice5_y_net,
    in_7 => slice6_y_net,
    in_8 => slice7_y_net,
    in_9 => slice8_y_net,
    in_10 => slice9_y_net,
    in_11 => slice10_y_net,
    in_12 => slice11_y_net,
    in_13 => slice12_y_net,
    in_14 => slice13_y_net,
    in_15 => slice14_y_net,
    in_16 => slice15_y_net,
    out_1 => reinterpret0_output_port_net,
    out_2 => reinterpret1_output_port_net,
    out_3 => reinterpret2_output_port_net,
    out_4 => reinterpret3_output_port_net,
    out_5 => reinterpret4_output_port_net,
    out_6 => reinterpret5_output_port_net,
    out_7 => reinterpret6_output_port_net,
    out_8 => reinterpret7_output_port_net,
    out_9 => reinterpret8_output_port_net,
    out_10 => reinterpret9_output_port_net,
    out_11 => reinterpret10_output_port_net,
    out_12 => reinterpret11_output_port_net,
    out_13 => reinterpret12_output_port_net,
    out_14 => reinterpret13_output_port_net,
    out_15 => reinterpret14_output_port_net,
    out_16 => reinterpret15_output_port_net
  );
  constant0 : entity xil_defaultlib.sysgen_constant_0714509e7f 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant0_op_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_31aefdfd97 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  constant2 : entity xil_defaultlib.sysgen_constant_de9059c03f 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant2_op_net
  );
  dpram_fir_coeffs_3 : entity xil_defaultlib.psb3_0_xltdpram 
  generic map (
    addr_width_b => 8,
    clocking_mode => "common_clock",
    data_width_b => 256,
    latency => 2,
    mem_init_file => "xpm_8f920b_vivado.mem",
    mem_size => 65536,
    mem_type => "block",
    read_reset_a => "0",
    read_reset_b => "0",
    width => 256,
    width_addr => 8,
    write_mode_a => "no_change",
    write_mode_b => "no_change"
  )
  port map (
    ena => "1",
    enb => "1",
    rsta => "0",
    rstb => "0",
    addra => read_addr_op_net,
    dina => constant1_op_net,
    wea => constant2_op_net,
    addrb => constant0_op_net,
    dinb => constant1_op_net,
    web => constant2_op_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dpram_fir_coeffs_3_douta_net,
    doutb => dpram_fir_coeffs_3_doutb_net
  );
  read_addr : entity xil_defaultlib.psb3_0_xlcounter_free 
  generic map (
    core_name0 => "psb3_0_c_counter_binary_v12_0_i0",
    op_arith => xlUnsigned,
    op_width => 8
  )
  port map (
    clr => '0',
    rst => gin_tl_reset_net,
    en => delay8_q_net,
    clk => clk_net,
    ce => ce_net,
    op => read_addr_op_net
  );
end structural;
-- Generated from Simulink block PSB3_0/DPRAM_FIR_Coeffs_4/Scalar to Vector
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_scalar_to_vector_x2 is
  port (
    i : in std_logic_vector( 256-1 downto 0 );
    o_1 : out std_logic_vector( 16-1 downto 0 );
    o_2 : out std_logic_vector( 16-1 downto 0 );
    o_3 : out std_logic_vector( 16-1 downto 0 );
    o_4 : out std_logic_vector( 16-1 downto 0 );
    o_5 : out std_logic_vector( 16-1 downto 0 );
    o_6 : out std_logic_vector( 16-1 downto 0 );
    o_7 : out std_logic_vector( 16-1 downto 0 );
    o_8 : out std_logic_vector( 16-1 downto 0 );
    o_9 : out std_logic_vector( 16-1 downto 0 );
    o_10 : out std_logic_vector( 16-1 downto 0 );
    o_11 : out std_logic_vector( 16-1 downto 0 );
    o_12 : out std_logic_vector( 16-1 downto 0 );
    o_13 : out std_logic_vector( 16-1 downto 0 );
    o_14 : out std_logic_vector( 16-1 downto 0 );
    o_15 : out std_logic_vector( 16-1 downto 0 );
    o_16 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_scalar_to_vector_x2;
architecture structural of psb3_0_scalar_to_vector_x2 is 
  signal slice0_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 16-1 downto 0 );
  signal dpram_fir_coeffs_4_douta_net : std_logic_vector( 256-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 16-1 downto 0 );
begin
  o_1 <= slice0_y_net;
  o_2 <= slice1_y_net;
  o_3 <= slice2_y_net;
  o_4 <= slice3_y_net;
  o_5 <= slice4_y_net;
  o_6 <= slice5_y_net;
  o_7 <= slice6_y_net;
  o_8 <= slice7_y_net;
  o_9 <= slice8_y_net;
  o_10 <= slice9_y_net;
  o_11 <= slice10_y_net;
  o_12 <= slice11_y_net;
  o_13 <= slice12_y_net;
  o_14 <= slice13_y_net;
  o_15 <= slice14_y_net;
  o_16 <= slice15_y_net;
  dpram_fir_coeffs_4_douta_net <= i;
  slice0 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 15,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => dpram_fir_coeffs_4_douta_net,
    y => slice0_y_net
  );
  slice1 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 16,
    new_msb => 31,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => dpram_fir_coeffs_4_douta_net,
    y => slice1_y_net
  );
  slice2 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 32,
    new_msb => 47,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => dpram_fir_coeffs_4_douta_net,
    y => slice2_y_net
  );
  slice3 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 48,
    new_msb => 63,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => dpram_fir_coeffs_4_douta_net,
    y => slice3_y_net
  );
  slice4 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 64,
    new_msb => 79,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => dpram_fir_coeffs_4_douta_net,
    y => slice4_y_net
  );
  slice5 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 80,
    new_msb => 95,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => dpram_fir_coeffs_4_douta_net,
    y => slice5_y_net
  );
  slice6 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 96,
    new_msb => 111,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => dpram_fir_coeffs_4_douta_net,
    y => slice6_y_net
  );
  slice7 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 112,
    new_msb => 127,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => dpram_fir_coeffs_4_douta_net,
    y => slice7_y_net
  );
  slice8 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 128,
    new_msb => 143,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => dpram_fir_coeffs_4_douta_net,
    y => slice8_y_net
  );
  slice9 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 144,
    new_msb => 159,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => dpram_fir_coeffs_4_douta_net,
    y => slice9_y_net
  );
  slice10 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 160,
    new_msb => 175,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => dpram_fir_coeffs_4_douta_net,
    y => slice10_y_net
  );
  slice11 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 176,
    new_msb => 191,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => dpram_fir_coeffs_4_douta_net,
    y => slice11_y_net
  );
  slice12 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 192,
    new_msb => 207,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => dpram_fir_coeffs_4_douta_net,
    y => slice12_y_net
  );
  slice13 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 208,
    new_msb => 223,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => dpram_fir_coeffs_4_douta_net,
    y => slice13_y_net
  );
  slice14 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 224,
    new_msb => 239,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => dpram_fir_coeffs_4_douta_net,
    y => slice14_y_net
  );
  slice15 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 240,
    new_msb => 255,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => dpram_fir_coeffs_4_douta_net,
    y => slice15_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/DPRAM_FIR_Coeffs_4/Vector Reinterpret
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_reinterpret_x2 is
  port (
    in_1 : in std_logic_vector( 16-1 downto 0 );
    in_2 : in std_logic_vector( 16-1 downto 0 );
    in_3 : in std_logic_vector( 16-1 downto 0 );
    in_4 : in std_logic_vector( 16-1 downto 0 );
    in_5 : in std_logic_vector( 16-1 downto 0 );
    in_6 : in std_logic_vector( 16-1 downto 0 );
    in_7 : in std_logic_vector( 16-1 downto 0 );
    in_8 : in std_logic_vector( 16-1 downto 0 );
    in_9 : in std_logic_vector( 16-1 downto 0 );
    in_10 : in std_logic_vector( 16-1 downto 0 );
    in_11 : in std_logic_vector( 16-1 downto 0 );
    in_12 : in std_logic_vector( 16-1 downto 0 );
    in_13 : in std_logic_vector( 16-1 downto 0 );
    in_14 : in std_logic_vector( 16-1 downto 0 );
    in_15 : in std_logic_vector( 16-1 downto 0 );
    in_16 : in std_logic_vector( 16-1 downto 0 );
    out_1 : out std_logic_vector( 16-1 downto 0 );
    out_2 : out std_logic_vector( 16-1 downto 0 );
    out_3 : out std_logic_vector( 16-1 downto 0 );
    out_4 : out std_logic_vector( 16-1 downto 0 );
    out_5 : out std_logic_vector( 16-1 downto 0 );
    out_6 : out std_logic_vector( 16-1 downto 0 );
    out_7 : out std_logic_vector( 16-1 downto 0 );
    out_8 : out std_logic_vector( 16-1 downto 0 );
    out_9 : out std_logic_vector( 16-1 downto 0 );
    out_10 : out std_logic_vector( 16-1 downto 0 );
    out_11 : out std_logic_vector( 16-1 downto 0 );
    out_12 : out std_logic_vector( 16-1 downto 0 );
    out_13 : out std_logic_vector( 16-1 downto 0 );
    out_14 : out std_logic_vector( 16-1 downto 0 );
    out_15 : out std_logic_vector( 16-1 downto 0 );
    out_16 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_vector_reinterpret_x2;
architecture structural of psb3_0_vector_reinterpret_x2 is 
  signal slice7_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 16-1 downto 0 );
begin
  out_1 <= reinterpret0_output_port_net;
  out_2 <= reinterpret1_output_port_net;
  out_3 <= reinterpret2_output_port_net;
  out_4 <= reinterpret3_output_port_net;
  out_5 <= reinterpret4_output_port_net;
  out_6 <= reinterpret5_output_port_net;
  out_7 <= reinterpret6_output_port_net;
  out_8 <= reinterpret7_output_port_net;
  out_9 <= reinterpret8_output_port_net;
  out_10 <= reinterpret9_output_port_net;
  out_11 <= reinterpret10_output_port_net;
  out_12 <= reinterpret11_output_port_net;
  out_13 <= reinterpret12_output_port_net;
  out_14 <= reinterpret13_output_port_net;
  out_15 <= reinterpret14_output_port_net;
  out_16 <= reinterpret15_output_port_net;
  slice0_y_net <= in_1;
  slice1_y_net <= in_2;
  slice2_y_net <= in_3;
  slice3_y_net <= in_4;
  slice4_y_net <= in_5;
  slice5_y_net <= in_6;
  slice6_y_net <= in_7;
  slice7_y_net <= in_8;
  slice8_y_net <= in_9;
  slice9_y_net <= in_10;
  slice10_y_net <= in_11;
  slice11_y_net <= in_12;
  slice12_y_net <= in_13;
  slice13_y_net <= in_14;
  slice14_y_net <= in_15;
  slice15_y_net <= in_16;
  reinterpret0 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice0_y_net,
    output_port => reinterpret0_output_port_net
  );
  reinterpret1 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice1_y_net,
    output_port => reinterpret1_output_port_net
  );
  reinterpret2 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice2_y_net,
    output_port => reinterpret2_output_port_net
  );
  reinterpret3 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice3_y_net,
    output_port => reinterpret3_output_port_net
  );
  reinterpret4 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice4_y_net,
    output_port => reinterpret4_output_port_net
  );
  reinterpret5 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice5_y_net,
    output_port => reinterpret5_output_port_net
  );
  reinterpret6 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice6_y_net,
    output_port => reinterpret6_output_port_net
  );
  reinterpret7 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice7_y_net,
    output_port => reinterpret7_output_port_net
  );
  reinterpret8 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice8_y_net,
    output_port => reinterpret8_output_port_net
  );
  reinterpret9 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice9_y_net,
    output_port => reinterpret9_output_port_net
  );
  reinterpret10 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice10_y_net,
    output_port => reinterpret10_output_port_net
  );
  reinterpret11 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice11_y_net,
    output_port => reinterpret11_output_port_net
  );
  reinterpret12 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice12_y_net,
    output_port => reinterpret12_output_port_net
  );
  reinterpret13 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice13_y_net,
    output_port => reinterpret13_output_port_net
  );
  reinterpret14 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice14_y_net,
    output_port => reinterpret14_output_port_net
  );
  reinterpret15 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice15_y_net,
    output_port => reinterpret15_output_port_net
  );
end structural;
-- Generated from Simulink block PSB3_0/DPRAM_FIR_Coeffs_4
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_dpram_fir_coeffs_4 is
  port (
    in_rst : in std_logic_vector( 1-1 downto 0 );
    in_en : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    out_fir_coeffs_1 : out std_logic_vector( 16-1 downto 0 );
    out_fir_coeffs_2 : out std_logic_vector( 16-1 downto 0 );
    out_fir_coeffs_3 : out std_logic_vector( 16-1 downto 0 );
    out_fir_coeffs_4 : out std_logic_vector( 16-1 downto 0 );
    out_fir_coeffs_5 : out std_logic_vector( 16-1 downto 0 );
    out_fir_coeffs_6 : out std_logic_vector( 16-1 downto 0 );
    out_fir_coeffs_7 : out std_logic_vector( 16-1 downto 0 );
    out_fir_coeffs_8 : out std_logic_vector( 16-1 downto 0 );
    out_fir_coeffs_9 : out std_logic_vector( 16-1 downto 0 );
    out_fir_coeffs_10 : out std_logic_vector( 16-1 downto 0 );
    out_fir_coeffs_11 : out std_logic_vector( 16-1 downto 0 );
    out_fir_coeffs_12 : out std_logic_vector( 16-1 downto 0 );
    out_fir_coeffs_13 : out std_logic_vector( 16-1 downto 0 );
    out_fir_coeffs_14 : out std_logic_vector( 16-1 downto 0 );
    out_fir_coeffs_15 : out std_logic_vector( 16-1 downto 0 );
    out_fir_coeffs_16 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_dpram_fir_coeffs_4;
architecture structural of psb3_0_dpram_fir_coeffs_4 is 
  signal ce_net : std_logic;
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal gin_tl_reset_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 16-1 downto 0 );
  signal clk_net : std_logic;
  signal slice6_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 16-1 downto 0 );
  signal dpram_fir_coeffs_4_douta_net : std_logic_vector( 256-1 downto 0 );
  signal constant0_op_net : std_logic_vector( 8-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 256-1 downto 0 );
  signal constant2_op_net : std_logic_vector( 1-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 16-1 downto 0 );
  signal dpram_fir_coeffs_4_doutb_net : std_logic_vector( 256-1 downto 0 );
  signal read_addr_op_net : std_logic_vector( 8-1 downto 0 );
begin
  out_fir_coeffs_1 <= reinterpret0_output_port_net;
  out_fir_coeffs_2 <= reinterpret1_output_port_net;
  out_fir_coeffs_3 <= reinterpret2_output_port_net;
  out_fir_coeffs_4 <= reinterpret3_output_port_net;
  out_fir_coeffs_5 <= reinterpret4_output_port_net;
  out_fir_coeffs_6 <= reinterpret5_output_port_net;
  out_fir_coeffs_7 <= reinterpret6_output_port_net;
  out_fir_coeffs_8 <= reinterpret7_output_port_net;
  out_fir_coeffs_9 <= reinterpret8_output_port_net;
  out_fir_coeffs_10 <= reinterpret9_output_port_net;
  out_fir_coeffs_11 <= reinterpret10_output_port_net;
  out_fir_coeffs_12 <= reinterpret11_output_port_net;
  out_fir_coeffs_13 <= reinterpret12_output_port_net;
  out_fir_coeffs_14 <= reinterpret13_output_port_net;
  out_fir_coeffs_15 <= reinterpret14_output_port_net;
  out_fir_coeffs_16 <= reinterpret15_output_port_net;
  gin_tl_reset_net <= in_rst;
  delay8_q_net <= in_en;
  clk_net <= clk_1;
  ce_net <= ce_1;
  scalar_to_vector : entity xil_defaultlib.psb3_0_scalar_to_vector_x2 
  port map (
    i => dpram_fir_coeffs_4_douta_net,
    o_1 => slice0_y_net,
    o_2 => slice1_y_net,
    o_3 => slice2_y_net,
    o_4 => slice3_y_net,
    o_5 => slice4_y_net,
    o_6 => slice5_y_net,
    o_7 => slice6_y_net,
    o_8 => slice7_y_net,
    o_9 => slice8_y_net,
    o_10 => slice9_y_net,
    o_11 => slice10_y_net,
    o_12 => slice11_y_net,
    o_13 => slice12_y_net,
    o_14 => slice13_y_net,
    o_15 => slice14_y_net,
    o_16 => slice15_y_net
  );
  vector_reinterpret : entity xil_defaultlib.psb3_0_vector_reinterpret_x2 
  port map (
    in_1 => slice0_y_net,
    in_2 => slice1_y_net,
    in_3 => slice2_y_net,
    in_4 => slice3_y_net,
    in_5 => slice4_y_net,
    in_6 => slice5_y_net,
    in_7 => slice6_y_net,
    in_8 => slice7_y_net,
    in_9 => slice8_y_net,
    in_10 => slice9_y_net,
    in_11 => slice10_y_net,
    in_12 => slice11_y_net,
    in_13 => slice12_y_net,
    in_14 => slice13_y_net,
    in_15 => slice14_y_net,
    in_16 => slice15_y_net,
    out_1 => reinterpret0_output_port_net,
    out_2 => reinterpret1_output_port_net,
    out_3 => reinterpret2_output_port_net,
    out_4 => reinterpret3_output_port_net,
    out_5 => reinterpret4_output_port_net,
    out_6 => reinterpret5_output_port_net,
    out_7 => reinterpret6_output_port_net,
    out_8 => reinterpret7_output_port_net,
    out_9 => reinterpret8_output_port_net,
    out_10 => reinterpret9_output_port_net,
    out_11 => reinterpret10_output_port_net,
    out_12 => reinterpret11_output_port_net,
    out_13 => reinterpret12_output_port_net,
    out_14 => reinterpret13_output_port_net,
    out_15 => reinterpret14_output_port_net,
    out_16 => reinterpret15_output_port_net
  );
  constant0 : entity xil_defaultlib.sysgen_constant_0714509e7f 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant0_op_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_31aefdfd97 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  constant2 : entity xil_defaultlib.sysgen_constant_de9059c03f 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant2_op_net
  );
  dpram_fir_coeffs_4 : entity xil_defaultlib.psb3_0_xltdpram 
  generic map (
    addr_width_b => 8,
    clocking_mode => "common_clock",
    data_width_b => 256,
    latency => 2,
    mem_init_file => "xpm_912a53_vivado.mem",
    mem_size => 65536,
    mem_type => "block",
    read_reset_a => "0",
    read_reset_b => "0",
    width => 256,
    width_addr => 8,
    write_mode_a => "no_change",
    write_mode_b => "no_change"
  )
  port map (
    ena => "1",
    enb => "1",
    rsta => "0",
    rstb => "0",
    addra => read_addr_op_net,
    dina => constant1_op_net,
    wea => constant2_op_net,
    addrb => constant0_op_net,
    dinb => constant1_op_net,
    web => constant2_op_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dpram_fir_coeffs_4_douta_net,
    doutb => dpram_fir_coeffs_4_doutb_net
  );
  read_addr : entity xil_defaultlib.psb3_0_xlcounter_free 
  generic map (
    core_name0 => "psb3_0_c_counter_binary_v12_0_i0",
    op_arith => xlUnsigned,
    op_width => 8
  )
  port map (
    clr => '0',
    rst => gin_tl_reset_net,
    en => delay8_q_net,
    clk => clk_net,
    ce => ce_net,
    op => read_addr_op_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Overflow Detector add_im_1/Vector Delay
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_delay is
  port (
    d_1 : in std_logic_vector( 1-1 downto 0 );
    d_2 : in std_logic_vector( 1-1 downto 0 );
    d_3 : in std_logic_vector( 1-1 downto 0 );
    d_4 : in std_logic_vector( 1-1 downto 0 );
    d_5 : in std_logic_vector( 1-1 downto 0 );
    d_6 : in std_logic_vector( 1-1 downto 0 );
    d_7 : in std_logic_vector( 1-1 downto 0 );
    d_8 : in std_logic_vector( 1-1 downto 0 );
    d_9 : in std_logic_vector( 1-1 downto 0 );
    d_10 : in std_logic_vector( 1-1 downto 0 );
    d_11 : in std_logic_vector( 1-1 downto 0 );
    d_12 : in std_logic_vector( 1-1 downto 0 );
    d_13 : in std_logic_vector( 1-1 downto 0 );
    d_14 : in std_logic_vector( 1-1 downto 0 );
    d_15 : in std_logic_vector( 1-1 downto 0 );
    d_16 : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    q_1 : out std_logic_vector( 1-1 downto 0 );
    q_2 : out std_logic_vector( 1-1 downto 0 );
    q_3 : out std_logic_vector( 1-1 downto 0 );
    q_4 : out std_logic_vector( 1-1 downto 0 );
    q_5 : out std_logic_vector( 1-1 downto 0 );
    q_6 : out std_logic_vector( 1-1 downto 0 );
    q_7 : out std_logic_vector( 1-1 downto 0 );
    q_8 : out std_logic_vector( 1-1 downto 0 );
    q_9 : out std_logic_vector( 1-1 downto 0 );
    q_10 : out std_logic_vector( 1-1 downto 0 );
    q_11 : out std_logic_vector( 1-1 downto 0 );
    q_12 : out std_logic_vector( 1-1 downto 0 );
    q_13 : out std_logic_vector( 1-1 downto 0 );
    q_14 : out std_logic_vector( 1-1 downto 0 );
    q_15 : out std_logic_vector( 1-1 downto 0 );
    q_16 : out std_logic_vector( 1-1 downto 0 )
  );
end psb3_0_vector_delay;
architecture structural of psb3_0_vector_delay is 
  signal delay5_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay9_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay11_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay13_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay0_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay7_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay14_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay15_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay10_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay12_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal ce_net : std_logic;
begin
  q_1 <= delay0_q_net;
  q_2 <= delay1_q_net;
  q_3 <= delay2_q_net;
  q_4 <= delay3_q_net;
  q_5 <= delay4_q_net;
  q_6 <= delay5_q_net;
  q_7 <= delay6_q_net;
  q_8 <= delay7_q_net;
  q_9 <= delay8_q_net;
  q_10 <= delay9_q_net;
  q_11 <= delay10_q_net;
  q_12 <= delay11_q_net;
  q_13 <= delay12_q_net;
  q_14 <= delay13_q_net;
  q_15 <= delay14_q_net;
  q_16 <= delay15_q_net;
  slice0_y_net <= d_1;
  slice1_y_net <= d_2;
  slice2_y_net <= d_3;
  slice3_y_net <= d_4;
  slice4_y_net <= d_5;
  slice5_y_net <= d_6;
  slice6_y_net <= d_7;
  slice7_y_net <= d_8;
  slice8_y_net <= d_9;
  slice9_y_net <= d_10;
  slice10_y_net <= d_11;
  slice11_y_net <= d_12;
  slice12_y_net <= d_13;
  slice13_y_net <= d_14;
  slice14_y_net <= d_15;
  slice15_y_net <= d_16;
  clk_net <= clk_1;
  ce_net <= ce_1;
  delay0 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice0_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay0_q_net
  );
  delay1 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice2_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay3 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice3_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  delay4 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice4_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net
  );
  delay5 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice5_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  delay6 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice6_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay6_q_net
  );
  delay7 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice7_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay7_q_net
  );
  delay8 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice8_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay8_q_net
  );
  delay9 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice9_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay9_q_net
  );
  delay10 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice10_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay10_q_net
  );
  delay11 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice11_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay11_q_net
  );
  delay12 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice12_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay12_q_net
  );
  delay13 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice13_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay13_q_net
  );
  delay14 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice14_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay14_q_net
  );
  delay15 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice15_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay15_q_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Overflow Detector add_im_1/Vector Delay1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_delay1 is
  port (
    d_1 : in std_logic_vector( 1-1 downto 0 );
    d_2 : in std_logic_vector( 1-1 downto 0 );
    d_3 : in std_logic_vector( 1-1 downto 0 );
    d_4 : in std_logic_vector( 1-1 downto 0 );
    d_5 : in std_logic_vector( 1-1 downto 0 );
    d_6 : in std_logic_vector( 1-1 downto 0 );
    d_7 : in std_logic_vector( 1-1 downto 0 );
    d_8 : in std_logic_vector( 1-1 downto 0 );
    d_9 : in std_logic_vector( 1-1 downto 0 );
    d_10 : in std_logic_vector( 1-1 downto 0 );
    d_11 : in std_logic_vector( 1-1 downto 0 );
    d_12 : in std_logic_vector( 1-1 downto 0 );
    d_13 : in std_logic_vector( 1-1 downto 0 );
    d_14 : in std_logic_vector( 1-1 downto 0 );
    d_15 : in std_logic_vector( 1-1 downto 0 );
    d_16 : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    q_1 : out std_logic_vector( 1-1 downto 0 );
    q_2 : out std_logic_vector( 1-1 downto 0 );
    q_3 : out std_logic_vector( 1-1 downto 0 );
    q_4 : out std_logic_vector( 1-1 downto 0 );
    q_5 : out std_logic_vector( 1-1 downto 0 );
    q_6 : out std_logic_vector( 1-1 downto 0 );
    q_7 : out std_logic_vector( 1-1 downto 0 );
    q_8 : out std_logic_vector( 1-1 downto 0 );
    q_9 : out std_logic_vector( 1-1 downto 0 );
    q_10 : out std_logic_vector( 1-1 downto 0 );
    q_11 : out std_logic_vector( 1-1 downto 0 );
    q_12 : out std_logic_vector( 1-1 downto 0 );
    q_13 : out std_logic_vector( 1-1 downto 0 );
    q_14 : out std_logic_vector( 1-1 downto 0 );
    q_15 : out std_logic_vector( 1-1 downto 0 );
    q_16 : out std_logic_vector( 1-1 downto 0 )
  );
end psb3_0_vector_delay1;
architecture structural of psb3_0_vector_delay1 is 
  signal slice6_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay0_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay15_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay11_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay13_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay14_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay12_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay7_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay9_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay10_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal slice14_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
begin
  q_1 <= delay0_q_net;
  q_2 <= delay1_q_net;
  q_3 <= delay2_q_net;
  q_4 <= delay3_q_net;
  q_5 <= delay4_q_net;
  q_6 <= delay5_q_net;
  q_7 <= delay6_q_net;
  q_8 <= delay7_q_net;
  q_9 <= delay8_q_net;
  q_10 <= delay9_q_net;
  q_11 <= delay10_q_net;
  q_12 <= delay11_q_net;
  q_13 <= delay12_q_net;
  q_14 <= delay13_q_net;
  q_15 <= delay14_q_net;
  q_16 <= delay15_q_net;
  slice0_y_net <= d_1;
  slice1_y_net <= d_2;
  slice2_y_net <= d_3;
  slice3_y_net <= d_4;
  slice4_y_net <= d_5;
  slice5_y_net <= d_6;
  slice6_y_net <= d_7;
  slice7_y_net <= d_8;
  slice8_y_net <= d_9;
  slice9_y_net <= d_10;
  slice10_y_net <= d_11;
  slice11_y_net <= d_12;
  slice12_y_net <= d_13;
  slice13_y_net <= d_14;
  slice14_y_net <= d_15;
  slice15_y_net <= d_16;
  clk_net <= clk_1;
  ce_net <= ce_1;
  delay0 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice0_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay0_q_net
  );
  delay1 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice2_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay3 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice3_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  delay4 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice4_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net
  );
  delay5 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice5_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  delay6 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice6_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay6_q_net
  );
  delay7 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice7_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay7_q_net
  );
  delay8 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice8_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay8_q_net
  );
  delay9 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice9_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay9_q_net
  );
  delay10 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice10_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay10_q_net
  );
  delay11 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice11_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay11_q_net
  );
  delay12 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice12_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay12_q_net
  );
  delay13 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice13_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay13_q_net
  );
  delay14 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice14_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay14_q_net
  );
  delay15 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice15_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay15_q_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Overflow Detector add_im_1/Vector Slice
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_slice is
  port (
    in_1 : in std_logic_vector( 16-1 downto 0 );
    in_2 : in std_logic_vector( 16-1 downto 0 );
    in_3 : in std_logic_vector( 16-1 downto 0 );
    in_4 : in std_logic_vector( 16-1 downto 0 );
    in_5 : in std_logic_vector( 16-1 downto 0 );
    in_6 : in std_logic_vector( 16-1 downto 0 );
    in_7 : in std_logic_vector( 16-1 downto 0 );
    in_8 : in std_logic_vector( 16-1 downto 0 );
    in_9 : in std_logic_vector( 16-1 downto 0 );
    in_10 : in std_logic_vector( 16-1 downto 0 );
    in_11 : in std_logic_vector( 16-1 downto 0 );
    in_12 : in std_logic_vector( 16-1 downto 0 );
    in_13 : in std_logic_vector( 16-1 downto 0 );
    in_14 : in std_logic_vector( 16-1 downto 0 );
    in_15 : in std_logic_vector( 16-1 downto 0 );
    in_16 : in std_logic_vector( 16-1 downto 0 );
    out_1 : out std_logic_vector( 1-1 downto 0 );
    out_2 : out std_logic_vector( 1-1 downto 0 );
    out_3 : out std_logic_vector( 1-1 downto 0 );
    out_4 : out std_logic_vector( 1-1 downto 0 );
    out_5 : out std_logic_vector( 1-1 downto 0 );
    out_6 : out std_logic_vector( 1-1 downto 0 );
    out_7 : out std_logic_vector( 1-1 downto 0 );
    out_8 : out std_logic_vector( 1-1 downto 0 );
    out_9 : out std_logic_vector( 1-1 downto 0 );
    out_10 : out std_logic_vector( 1-1 downto 0 );
    out_11 : out std_logic_vector( 1-1 downto 0 );
    out_12 : out std_logic_vector( 1-1 downto 0 );
    out_13 : out std_logic_vector( 1-1 downto 0 );
    out_14 : out std_logic_vector( 1-1 downto 0 );
    out_15 : out std_logic_vector( 1-1 downto 0 );
    out_16 : out std_logic_vector( 1-1 downto 0 )
  );
end psb3_0_vector_slice;
architecture structural of psb3_0_vector_slice is 
  signal slice5_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 1-1 downto 0 );
  signal mult5_p_net : std_logic_vector( 16-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 1-1 downto 0 );
  signal mult4_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult12_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult8_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult7_p_net : std_logic_vector( 16-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 1-1 downto 0 );
  signal mult2_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult1_p_net : std_logic_vector( 16-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 1-1 downto 0 );
  signal mult14_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult6_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult10_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult11_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult3_p_net : std_logic_vector( 16-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 1-1 downto 0 );
  signal mult9_p_net : std_logic_vector( 16-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 1-1 downto 0 );
  signal mult13_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult0_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult15_p_net : std_logic_vector( 16-1 downto 0 );
begin
  out_1 <= slice0_y_net;
  out_2 <= slice1_y_net;
  out_3 <= slice2_y_net;
  out_4 <= slice3_y_net;
  out_5 <= slice4_y_net;
  out_6 <= slice5_y_net;
  out_7 <= slice6_y_net;
  out_8 <= slice7_y_net;
  out_9 <= slice8_y_net;
  out_10 <= slice9_y_net;
  out_11 <= slice10_y_net;
  out_12 <= slice11_y_net;
  out_13 <= slice12_y_net;
  out_14 <= slice13_y_net;
  out_15 <= slice14_y_net;
  out_16 <= slice15_y_net;
  mult0_p_net <= in_1;
  mult1_p_net <= in_2;
  mult2_p_net <= in_3;
  mult3_p_net <= in_4;
  mult4_p_net <= in_5;
  mult5_p_net <= in_6;
  mult6_p_net <= in_7;
  mult7_p_net <= in_8;
  mult8_p_net <= in_9;
  mult9_p_net <= in_10;
  mult10_p_net <= in_11;
  mult11_p_net <= in_12;
  mult12_p_net <= in_13;
  mult13_p_net <= in_14;
  mult14_p_net <= in_15;
  mult15_p_net <= in_16;
  slice0 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult0_p_net,
    y => slice0_y_net
  );
  slice1 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult1_p_net,
    y => slice1_y_net
  );
  slice2 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult2_p_net,
    y => slice2_y_net
  );
  slice3 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult3_p_net,
    y => slice3_y_net
  );
  slice4 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult4_p_net,
    y => slice4_y_net
  );
  slice5 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult5_p_net,
    y => slice5_y_net
  );
  slice6 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult6_p_net,
    y => slice6_y_net
  );
  slice7 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult7_p_net,
    y => slice7_y_net
  );
  slice8 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult8_p_net,
    y => slice8_y_net
  );
  slice9 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult9_p_net,
    y => slice9_y_net
  );
  slice10 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult10_p_net,
    y => slice10_y_net
  );
  slice11 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult11_p_net,
    y => slice11_y_net
  );
  slice12 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult12_p_net,
    y => slice12_y_net
  );
  slice13 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult13_p_net,
    y => slice13_y_net
  );
  slice14 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult14_p_net,
    y => slice14_y_net
  );
  slice15 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult15_p_net,
    y => slice15_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Overflow Detector add_im_1/Vector Slice1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_slice1 is
  port (
    in_1 : in std_logic_vector( 16-1 downto 0 );
    in_2 : in std_logic_vector( 16-1 downto 0 );
    in_3 : in std_logic_vector( 16-1 downto 0 );
    in_4 : in std_logic_vector( 16-1 downto 0 );
    in_5 : in std_logic_vector( 16-1 downto 0 );
    in_6 : in std_logic_vector( 16-1 downto 0 );
    in_7 : in std_logic_vector( 16-1 downto 0 );
    in_8 : in std_logic_vector( 16-1 downto 0 );
    in_9 : in std_logic_vector( 16-1 downto 0 );
    in_10 : in std_logic_vector( 16-1 downto 0 );
    in_11 : in std_logic_vector( 16-1 downto 0 );
    in_12 : in std_logic_vector( 16-1 downto 0 );
    in_13 : in std_logic_vector( 16-1 downto 0 );
    in_14 : in std_logic_vector( 16-1 downto 0 );
    in_15 : in std_logic_vector( 16-1 downto 0 );
    in_16 : in std_logic_vector( 16-1 downto 0 );
    out_1 : out std_logic_vector( 1-1 downto 0 );
    out_2 : out std_logic_vector( 1-1 downto 0 );
    out_3 : out std_logic_vector( 1-1 downto 0 );
    out_4 : out std_logic_vector( 1-1 downto 0 );
    out_5 : out std_logic_vector( 1-1 downto 0 );
    out_6 : out std_logic_vector( 1-1 downto 0 );
    out_7 : out std_logic_vector( 1-1 downto 0 );
    out_8 : out std_logic_vector( 1-1 downto 0 );
    out_9 : out std_logic_vector( 1-1 downto 0 );
    out_10 : out std_logic_vector( 1-1 downto 0 );
    out_11 : out std_logic_vector( 1-1 downto 0 );
    out_12 : out std_logic_vector( 1-1 downto 0 );
    out_13 : out std_logic_vector( 1-1 downto 0 );
    out_14 : out std_logic_vector( 1-1 downto 0 );
    out_15 : out std_logic_vector( 1-1 downto 0 );
    out_16 : out std_logic_vector( 1-1 downto 0 )
  );
end psb3_0_vector_slice1;
architecture structural of psb3_0_vector_slice1 is 
  signal slice3_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
begin
  out_1 <= slice0_y_net;
  out_2 <= slice1_y_net;
  out_3 <= slice2_y_net;
  out_4 <= slice3_y_net;
  out_5 <= slice4_y_net;
  out_6 <= slice5_y_net;
  out_7 <= slice6_y_net;
  out_8 <= slice7_y_net;
  out_9 <= slice8_y_net;
  out_10 <= slice9_y_net;
  out_11 <= slice10_y_net;
  out_12 <= slice11_y_net;
  out_13 <= slice12_y_net;
  out_14 <= slice13_y_net;
  out_15 <= slice14_y_net;
  out_16 <= slice15_y_net;
  reinterpret0_output_port_net <= in_1;
  reinterpret1_output_port_net <= in_2;
  reinterpret2_output_port_net <= in_3;
  reinterpret3_output_port_net <= in_4;
  reinterpret4_output_port_net <= in_5;
  reinterpret5_output_port_net <= in_6;
  reinterpret6_output_port_net <= in_7;
  reinterpret7_output_port_net <= in_8;
  reinterpret8_output_port_net <= in_9;
  reinterpret9_output_port_net <= in_10;
  reinterpret10_output_port_net <= in_11;
  reinterpret11_output_port_net <= in_12;
  reinterpret12_output_port_net <= in_13;
  reinterpret13_output_port_net <= in_14;
  reinterpret14_output_port_net <= in_15;
  reinterpret15_output_port_net <= in_16;
  slice0 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret0_output_port_net,
    y => slice0_y_net
  );
  slice1 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret1_output_port_net,
    y => slice1_y_net
  );
  slice2 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret2_output_port_net,
    y => slice2_y_net
  );
  slice3 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret3_output_port_net,
    y => slice3_y_net
  );
  slice4 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret4_output_port_net,
    y => slice4_y_net
  );
  slice5 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret5_output_port_net,
    y => slice5_y_net
  );
  slice6 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret6_output_port_net,
    y => slice6_y_net
  );
  slice7 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret7_output_port_net,
    y => slice7_y_net
  );
  slice8 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret8_output_port_net,
    y => slice8_y_net
  );
  slice9 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret9_output_port_net,
    y => slice9_y_net
  );
  slice10 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret10_output_port_net,
    y => slice10_y_net
  );
  slice11 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret11_output_port_net,
    y => slice11_y_net
  );
  slice12 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret12_output_port_net,
    y => slice12_y_net
  );
  slice13 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret13_output_port_net,
    y => slice13_y_net
  );
  slice14 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret14_output_port_net,
    y => slice14_y_net
  );
  slice15 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret15_output_port_net,
    y => slice15_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Overflow Detector add_im_1/Vector Slice2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_slice2 is
  port (
    in_1 : in std_logic_vector( 16-1 downto 0 );
    in_2 : in std_logic_vector( 16-1 downto 0 );
    in_3 : in std_logic_vector( 16-1 downto 0 );
    in_4 : in std_logic_vector( 16-1 downto 0 );
    in_5 : in std_logic_vector( 16-1 downto 0 );
    in_6 : in std_logic_vector( 16-1 downto 0 );
    in_7 : in std_logic_vector( 16-1 downto 0 );
    in_8 : in std_logic_vector( 16-1 downto 0 );
    in_9 : in std_logic_vector( 16-1 downto 0 );
    in_10 : in std_logic_vector( 16-1 downto 0 );
    in_11 : in std_logic_vector( 16-1 downto 0 );
    in_12 : in std_logic_vector( 16-1 downto 0 );
    in_13 : in std_logic_vector( 16-1 downto 0 );
    in_14 : in std_logic_vector( 16-1 downto 0 );
    in_15 : in std_logic_vector( 16-1 downto 0 );
    in_16 : in std_logic_vector( 16-1 downto 0 );
    out_1 : out std_logic_vector( 1-1 downto 0 );
    out_2 : out std_logic_vector( 1-1 downto 0 );
    out_3 : out std_logic_vector( 1-1 downto 0 );
    out_4 : out std_logic_vector( 1-1 downto 0 );
    out_5 : out std_logic_vector( 1-1 downto 0 );
    out_6 : out std_logic_vector( 1-1 downto 0 );
    out_7 : out std_logic_vector( 1-1 downto 0 );
    out_8 : out std_logic_vector( 1-1 downto 0 );
    out_9 : out std_logic_vector( 1-1 downto 0 );
    out_10 : out std_logic_vector( 1-1 downto 0 );
    out_11 : out std_logic_vector( 1-1 downto 0 );
    out_12 : out std_logic_vector( 1-1 downto 0 );
    out_13 : out std_logic_vector( 1-1 downto 0 );
    out_14 : out std_logic_vector( 1-1 downto 0 );
    out_15 : out std_logic_vector( 1-1 downto 0 );
    out_16 : out std_logic_vector( 1-1 downto 0 )
  );
end psb3_0_vector_slice2;
architecture structural of psb3_0_vector_slice2 is 
  signal slice2_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 1-1 downto 0 );
  signal addsub11_s_net : std_logic_vector( 16-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 1-1 downto 0 );
  signal addsub10_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub12_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub13_s_net : std_logic_vector( 16-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 1-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 16-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 1-1 downto 0 );
  signal addsub5_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub7_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub8_s_net : std_logic_vector( 16-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 1-1 downto 0 );
  signal addsub9_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub3_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub14_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub0_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub15_s_net : std_logic_vector( 16-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 1-1 downto 0 );
  signal addsub6_s_net : std_logic_vector( 16-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 1-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 16-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 1-1 downto 0 );
begin
  out_1 <= slice0_y_net;
  out_2 <= slice1_y_net;
  out_3 <= slice2_y_net;
  out_4 <= slice3_y_net;
  out_5 <= slice4_y_net;
  out_6 <= slice5_y_net;
  out_7 <= slice6_y_net;
  out_8 <= slice7_y_net;
  out_9 <= slice8_y_net;
  out_10 <= slice9_y_net;
  out_11 <= slice10_y_net;
  out_12 <= slice11_y_net;
  out_13 <= slice12_y_net;
  out_14 <= slice13_y_net;
  out_15 <= slice14_y_net;
  out_16 <= slice15_y_net;
  addsub0_s_net <= in_1;
  addsub1_s_net <= in_2;
  addsub2_s_net <= in_3;
  addsub3_s_net <= in_4;
  addsub4_s_net <= in_5;
  addsub5_s_net <= in_6;
  addsub6_s_net <= in_7;
  addsub7_s_net <= in_8;
  addsub8_s_net <= in_9;
  addsub9_s_net <= in_10;
  addsub10_s_net <= in_11;
  addsub11_s_net <= in_12;
  addsub12_s_net <= in_13;
  addsub13_s_net <= in_14;
  addsub14_s_net <= in_15;
  addsub15_s_net <= in_16;
  slice0 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub0_s_net,
    y => slice0_y_net
  );
  slice1 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub1_s_net,
    y => slice1_y_net
  );
  slice2 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub2_s_net,
    y => slice2_y_net
  );
  slice3 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub3_s_net,
    y => slice3_y_net
  );
  slice4 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub4_s_net,
    y => slice4_y_net
  );
  slice5 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub5_s_net,
    y => slice5_y_net
  );
  slice6 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub6_s_net,
    y => slice6_y_net
  );
  slice7 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub7_s_net,
    y => slice7_y_net
  );
  slice8 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub8_s_net,
    y => slice8_y_net
  );
  slice9 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub9_s_net,
    y => slice9_y_net
  );
  slice10 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub10_s_net,
    y => slice10_y_net
  );
  slice11 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub11_s_net,
    y => slice11_y_net
  );
  slice12 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub12_s_net,
    y => slice12_y_net
  );
  slice13 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub13_s_net,
    y => slice13_y_net
  );
  slice14 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub14_s_net,
    y => slice14_y_net
  );
  slice15 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub15_s_net,
    y => slice15_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Overflow Detector add_im_1/Vector to Scalar
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_to_scalar is
  port (
    i_1 : in std_logic_vector( 1-1 downto 0 );
    i_2 : in std_logic_vector( 1-1 downto 0 );
    i_3 : in std_logic_vector( 1-1 downto 0 );
    i_4 : in std_logic_vector( 1-1 downto 0 );
    i_5 : in std_logic_vector( 1-1 downto 0 );
    i_6 : in std_logic_vector( 1-1 downto 0 );
    i_7 : in std_logic_vector( 1-1 downto 0 );
    i_8 : in std_logic_vector( 1-1 downto 0 );
    i_9 : in std_logic_vector( 1-1 downto 0 );
    i_10 : in std_logic_vector( 1-1 downto 0 );
    i_11 : in std_logic_vector( 1-1 downto 0 );
    i_12 : in std_logic_vector( 1-1 downto 0 );
    i_13 : in std_logic_vector( 1-1 downto 0 );
    i_14 : in std_logic_vector( 1-1 downto 0 );
    i_15 : in std_logic_vector( 1-1 downto 0 );
    i_16 : in std_logic_vector( 1-1 downto 0 );
    o : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_vector_to_scalar;
architecture structural of psb3_0_vector_to_scalar is 
  signal delay3_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay7_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay10_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay11_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay9_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay12_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay15_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 1-1 downto 0 );
  signal concat1_y_net : std_logic_vector( 16-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay13_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay14_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay0_q_net : std_logic_vector( 1-1 downto 0 );
begin
  o <= concat1_y_net;
  delay0_q_net <= i_1;
  delay1_q_net <= i_2;
  delay2_q_net <= i_3;
  delay3_q_net <= i_4;
  delay4_q_net <= i_5;
  delay5_q_net <= i_6;
  delay6_q_net <= i_7;
  delay7_q_net <= i_8;
  delay8_q_net <= i_9;
  delay9_q_net <= i_10;
  delay10_q_net <= i_11;
  delay11_q_net <= i_12;
  delay12_q_net <= i_13;
  delay13_q_net <= i_14;
  delay14_q_net <= i_15;
  delay15_q_net <= i_16;
  concat1 : entity xil_defaultlib.sysgen_concat_d977c66e35 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => delay15_q_net,
    in1 => delay14_q_net,
    in2 => delay13_q_net,
    in3 => delay12_q_net,
    in4 => delay11_q_net,
    in5 => delay10_q_net,
    in6 => delay9_q_net,
    in7 => delay8_q_net,
    in8 => delay7_q_net,
    in9 => delay6_q_net,
    in10 => delay5_q_net,
    in11 => delay4_q_net,
    in12 => delay3_q_net,
    in13 => delay2_q_net,
    in14 => delay1_q_net,
    in15 => delay0_q_net,
    y => concat1_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Overflow Detector add_im_1/Vector to Scalar1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_to_scalar1 is
  port (
    i_1 : in std_logic_vector( 1-1 downto 0 );
    i_2 : in std_logic_vector( 1-1 downto 0 );
    i_3 : in std_logic_vector( 1-1 downto 0 );
    i_4 : in std_logic_vector( 1-1 downto 0 );
    i_5 : in std_logic_vector( 1-1 downto 0 );
    i_6 : in std_logic_vector( 1-1 downto 0 );
    i_7 : in std_logic_vector( 1-1 downto 0 );
    i_8 : in std_logic_vector( 1-1 downto 0 );
    i_9 : in std_logic_vector( 1-1 downto 0 );
    i_10 : in std_logic_vector( 1-1 downto 0 );
    i_11 : in std_logic_vector( 1-1 downto 0 );
    i_12 : in std_logic_vector( 1-1 downto 0 );
    i_13 : in std_logic_vector( 1-1 downto 0 );
    i_14 : in std_logic_vector( 1-1 downto 0 );
    i_15 : in std_logic_vector( 1-1 downto 0 );
    i_16 : in std_logic_vector( 1-1 downto 0 );
    o : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_vector_to_scalar1;
architecture structural of psb3_0_vector_to_scalar1 is 
  signal delay14_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay13_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay15_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay0_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay11_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay10_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay12_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay9_q_net : std_logic_vector( 1-1 downto 0 );
  signal concat1_y_net : std_logic_vector( 16-1 downto 0 );
  signal delay7_q_net : std_logic_vector( 1-1 downto 0 );
begin
  o <= concat1_y_net;
  delay0_q_net <= i_1;
  delay1_q_net <= i_2;
  delay2_q_net <= i_3;
  delay3_q_net <= i_4;
  delay4_q_net <= i_5;
  delay5_q_net <= i_6;
  delay6_q_net <= i_7;
  delay7_q_net <= i_8;
  delay8_q_net <= i_9;
  delay9_q_net <= i_10;
  delay10_q_net <= i_11;
  delay11_q_net <= i_12;
  delay12_q_net <= i_13;
  delay13_q_net <= i_14;
  delay14_q_net <= i_15;
  delay15_q_net <= i_16;
  concat1 : entity xil_defaultlib.sysgen_concat_d977c66e35 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => delay15_q_net,
    in1 => delay14_q_net,
    in2 => delay13_q_net,
    in3 => delay12_q_net,
    in4 => delay11_q_net,
    in5 => delay10_q_net,
    in6 => delay9_q_net,
    in7 => delay8_q_net,
    in8 => delay7_q_net,
    in9 => delay6_q_net,
    in10 => delay5_q_net,
    in11 => delay4_q_net,
    in12 => delay3_q_net,
    in13 => delay2_q_net,
    in14 => delay1_q_net,
    in15 => delay0_q_net,
    y => concat1_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Overflow Detector add_im_1/Vector to Scalar2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_to_scalar2_x0 is
  port (
    i_1 : in std_logic_vector( 1-1 downto 0 );
    i_2 : in std_logic_vector( 1-1 downto 0 );
    i_3 : in std_logic_vector( 1-1 downto 0 );
    i_4 : in std_logic_vector( 1-1 downto 0 );
    i_5 : in std_logic_vector( 1-1 downto 0 );
    i_6 : in std_logic_vector( 1-1 downto 0 );
    i_7 : in std_logic_vector( 1-1 downto 0 );
    i_8 : in std_logic_vector( 1-1 downto 0 );
    i_9 : in std_logic_vector( 1-1 downto 0 );
    i_10 : in std_logic_vector( 1-1 downto 0 );
    i_11 : in std_logic_vector( 1-1 downto 0 );
    i_12 : in std_logic_vector( 1-1 downto 0 );
    i_13 : in std_logic_vector( 1-1 downto 0 );
    i_14 : in std_logic_vector( 1-1 downto 0 );
    i_15 : in std_logic_vector( 1-1 downto 0 );
    i_16 : in std_logic_vector( 1-1 downto 0 );
    o : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_vector_to_scalar2_x0;
architecture structural of psb3_0_vector_to_scalar2_x0 is 
  signal slice15_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 1-1 downto 0 );
  signal concat1_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 1-1 downto 0 );
begin
  o <= concat1_y_net;
  slice0_y_net <= i_1;
  slice1_y_net <= i_2;
  slice2_y_net <= i_3;
  slice3_y_net <= i_4;
  slice4_y_net <= i_5;
  slice5_y_net <= i_6;
  slice6_y_net <= i_7;
  slice7_y_net <= i_8;
  slice8_y_net <= i_9;
  slice9_y_net <= i_10;
  slice10_y_net <= i_11;
  slice11_y_net <= i_12;
  slice12_y_net <= i_13;
  slice13_y_net <= i_14;
  slice14_y_net <= i_15;
  slice15_y_net <= i_16;
  concat1 : entity xil_defaultlib.sysgen_concat_d977c66e35 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => slice15_y_net,
    in1 => slice14_y_net,
    in2 => slice13_y_net,
    in3 => slice12_y_net,
    in4 => slice11_y_net,
    in5 => slice10_y_net,
    in6 => slice9_y_net,
    in7 => slice8_y_net,
    in8 => slice7_y_net,
    in9 => slice6_y_net,
    in10 => slice5_y_net,
    in11 => slice4_y_net,
    in12 => slice3_y_net,
    in13 => slice2_y_net,
    in14 => slice1_y_net,
    in15 => slice0_y_net,
    y => concat1_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Overflow Detector add_im_1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_overflow_detector_add_im_1 is
  port (
    rst : in std_logic_vector( 1-1 downto 0 );
    a_1 : in std_logic_vector( 16-1 downto 0 );
    b_1 : in std_logic_vector( 16-1 downto 0 );
    s_1 : in std_logic_vector( 16-1 downto 0 );
    a_2 : in std_logic_vector( 16-1 downto 0 );
    a_3 : in std_logic_vector( 16-1 downto 0 );
    a_4 : in std_logic_vector( 16-1 downto 0 );
    a_5 : in std_logic_vector( 16-1 downto 0 );
    a_6 : in std_logic_vector( 16-1 downto 0 );
    a_7 : in std_logic_vector( 16-1 downto 0 );
    a_8 : in std_logic_vector( 16-1 downto 0 );
    a_9 : in std_logic_vector( 16-1 downto 0 );
    a_10 : in std_logic_vector( 16-1 downto 0 );
    a_11 : in std_logic_vector( 16-1 downto 0 );
    a_12 : in std_logic_vector( 16-1 downto 0 );
    a_13 : in std_logic_vector( 16-1 downto 0 );
    a_14 : in std_logic_vector( 16-1 downto 0 );
    a_15 : in std_logic_vector( 16-1 downto 0 );
    a_16 : in std_logic_vector( 16-1 downto 0 );
    b_2 : in std_logic_vector( 16-1 downto 0 );
    b_3 : in std_logic_vector( 16-1 downto 0 );
    b_4 : in std_logic_vector( 16-1 downto 0 );
    b_5 : in std_logic_vector( 16-1 downto 0 );
    b_6 : in std_logic_vector( 16-1 downto 0 );
    b_7 : in std_logic_vector( 16-1 downto 0 );
    b_8 : in std_logic_vector( 16-1 downto 0 );
    b_9 : in std_logic_vector( 16-1 downto 0 );
    b_10 : in std_logic_vector( 16-1 downto 0 );
    b_11 : in std_logic_vector( 16-1 downto 0 );
    b_12 : in std_logic_vector( 16-1 downto 0 );
    b_13 : in std_logic_vector( 16-1 downto 0 );
    b_14 : in std_logic_vector( 16-1 downto 0 );
    b_15 : in std_logic_vector( 16-1 downto 0 );
    b_16 : in std_logic_vector( 16-1 downto 0 );
    s_2 : in std_logic_vector( 16-1 downto 0 );
    s_3 : in std_logic_vector( 16-1 downto 0 );
    s_4 : in std_logic_vector( 16-1 downto 0 );
    s_5 : in std_logic_vector( 16-1 downto 0 );
    s_6 : in std_logic_vector( 16-1 downto 0 );
    s_7 : in std_logic_vector( 16-1 downto 0 );
    s_8 : in std_logic_vector( 16-1 downto 0 );
    s_9 : in std_logic_vector( 16-1 downto 0 );
    s_10 : in std_logic_vector( 16-1 downto 0 );
    s_11 : in std_logic_vector( 16-1 downto 0 );
    s_12 : in std_logic_vector( 16-1 downto 0 );
    s_13 : in std_logic_vector( 16-1 downto 0 );
    s_14 : in std_logic_vector( 16-1 downto 0 );
    s_15 : in std_logic_vector( 16-1 downto 0 );
    s_16 : in std_logic_vector( 16-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    ov : out std_logic_vector( 1-1 downto 0 )
  );
end psb3_0_overflow_detector_add_im_1;
architecture structural of psb3_0_overflow_detector_add_im_1 is 
  signal register_q_net : std_logic_vector( 1-1 downto 0 );
  signal gin_tl_reset_net : std_logic_vector( 1-1 downto 0 );
  signal mult0_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult13_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult3_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mult7_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mult11_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult15_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mult1_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mult5_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mult12_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mult4_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult14_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub0_s_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mult6_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult2_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mult10_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mult8_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mult9_p_net : std_logic_vector( 16-1 downto 0 );
  signal addsub12_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub8_s_net : std_logic_vector( 16-1 downto 0 );
  signal delay7_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay14_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal addsub11_s_net : std_logic_vector( 16-1 downto 0 );
  signal slice0_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal addsub13_s_net : std_logic_vector( 16-1 downto 0 );
  signal clk_net : std_logic;
  signal delay11_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice4_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal delay15_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal addsub7_s_net : std_logic_vector( 16-1 downto 0 );
  signal delay2_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal addsub5_s_net : std_logic_vector( 16-1 downto 0 );
  signal delay6_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice1_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal addsub6_s_net : std_logic_vector( 16-1 downto 0 );
  signal delay9_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice6_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal slice8_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal slice12_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal slice13_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal slice11_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal addsub14_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub9_s_net : std_logic_vector( 16-1 downto 0 );
  signal slice14_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal slice3_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice2_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal slice9_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal delay12_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub10_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub15_s_net : std_logic_vector( 16-1 downto 0 );
  signal ce_net : std_logic;
  signal delay3_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay5_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay8_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay0_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub3_s_net : std_logic_vector( 16-1 downto 0 );
  signal delay4_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay10_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay13_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice5_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal slice7_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal slice10_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay7_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice9_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice8_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice4_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay11_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay0_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice5_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice12_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice1_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice13_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice14_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 1-1 downto 0 );
  signal concat1_y_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal concat1_y_net : std_logic_vector( 16-1 downto 0 );
  signal delay15_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice3_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay12_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice6_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 1-1 downto 0 );
  signal concat1_y_net_x1 : std_logic_vector( 16-1 downto 0 );
  signal constant17_op_net : std_logic_vector( 1-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice0_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 1-1 downto 0 );
  signal convert_dout_net : std_logic_vector( 1-1 downto 0 );
  signal delay10_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay9_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice11_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay14_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice15_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay13_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice7_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice15_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice10_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice2_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 1-1 downto 0 );
  signal expression_dout_net : std_logic_vector( 1-1 downto 0 );
begin
  ov <= register_q_net;
  gin_tl_reset_net <= rst;
  mult0_p_net <= a_1;
  reinterpret0_output_port_net <= b_1;
  addsub0_s_net <= s_1;
  mult1_p_net <= a_2;
  mult2_p_net <= a_3;
  mult3_p_net <= a_4;
  mult4_p_net <= a_5;
  mult5_p_net <= a_6;
  mult6_p_net <= a_7;
  mult7_p_net <= a_8;
  mult8_p_net <= a_9;
  mult9_p_net <= a_10;
  mult10_p_net <= a_11;
  mult11_p_net <= a_12;
  mult12_p_net <= a_13;
  mult13_p_net <= a_14;
  mult14_p_net <= a_15;
  mult15_p_net <= a_16;
  reinterpret1_output_port_net <= b_2;
  reinterpret2_output_port_net <= b_3;
  reinterpret3_output_port_net <= b_4;
  reinterpret4_output_port_net <= b_5;
  reinterpret5_output_port_net <= b_6;
  reinterpret6_output_port_net <= b_7;
  reinterpret7_output_port_net <= b_8;
  reinterpret8_output_port_net <= b_9;
  reinterpret9_output_port_net <= b_10;
  reinterpret10_output_port_net <= b_11;
  reinterpret11_output_port_net <= b_12;
  reinterpret12_output_port_net <= b_13;
  reinterpret13_output_port_net <= b_14;
  reinterpret14_output_port_net <= b_15;
  reinterpret15_output_port_net <= b_16;
  addsub1_s_net <= s_2;
  addsub2_s_net <= s_3;
  addsub3_s_net <= s_4;
  addsub4_s_net <= s_5;
  addsub5_s_net <= s_6;
  addsub6_s_net <= s_7;
  addsub7_s_net <= s_8;
  addsub8_s_net <= s_9;
  addsub9_s_net <= s_10;
  addsub10_s_net <= s_11;
  addsub11_s_net <= s_12;
  addsub12_s_net <= s_13;
  addsub13_s_net <= s_14;
  addsub14_s_net <= s_15;
  addsub15_s_net <= s_16;
  clk_net <= clk_1;
  ce_net <= ce_1;
  vector_delay : entity xil_defaultlib.psb3_0_vector_delay 
  port map (
    d_1 => slice0_y_net_x1,
    d_2 => slice1_y_net_x1,
    d_3 => slice2_y_net_x1,
    d_4 => slice3_y_net_x1,
    d_5 => slice4_y_net_x1,
    d_6 => slice5_y_net_x1,
    d_7 => slice6_y_net_x1,
    d_8 => slice7_y_net_x1,
    d_9 => slice8_y_net_x1,
    d_10 => slice9_y_net_x1,
    d_11 => slice10_y_net_x1,
    d_12 => slice11_y_net_x1,
    d_13 => slice12_y_net_x1,
    d_14 => slice13_y_net_x1,
    d_15 => slice14_y_net_x1,
    d_16 => slice15_y_net_x1,
    clk_1 => clk_net,
    ce_1 => ce_net,
    q_1 => delay0_q_net_x0,
    q_2 => delay1_q_net_x0,
    q_3 => delay2_q_net_x0,
    q_4 => delay3_q_net_x0,
    q_5 => delay4_q_net_x0,
    q_6 => delay5_q_net_x0,
    q_7 => delay6_q_net_x0,
    q_8 => delay7_q_net_x0,
    q_9 => delay8_q_net_x0,
    q_10 => delay9_q_net_x0,
    q_11 => delay10_q_net_x0,
    q_12 => delay11_q_net_x0,
    q_13 => delay12_q_net_x0,
    q_14 => delay13_q_net_x0,
    q_15 => delay14_q_net_x0,
    q_16 => delay15_q_net_x0
  );
  vector_delay1 : entity xil_defaultlib.psb3_0_vector_delay1 
  port map (
    d_1 => slice0_y_net_x0,
    d_2 => slice1_y_net_x0,
    d_3 => slice2_y_net_x0,
    d_4 => slice3_y_net_x0,
    d_5 => slice4_y_net_x0,
    d_6 => slice5_y_net_x0,
    d_7 => slice6_y_net_x0,
    d_8 => slice7_y_net_x0,
    d_9 => slice8_y_net_x0,
    d_10 => slice9_y_net_x0,
    d_11 => slice10_y_net_x0,
    d_12 => slice11_y_net_x0,
    d_13 => slice12_y_net_x0,
    d_14 => slice13_y_net_x0,
    d_15 => slice14_y_net_x0,
    d_16 => slice15_y_net_x0,
    clk_1 => clk_net,
    ce_1 => ce_net,
    q_1 => delay0_q_net,
    q_2 => delay1_q_net,
    q_3 => delay2_q_net,
    q_4 => delay3_q_net,
    q_5 => delay4_q_net,
    q_6 => delay5_q_net,
    q_7 => delay6_q_net,
    q_8 => delay7_q_net,
    q_9 => delay8_q_net,
    q_10 => delay9_q_net,
    q_11 => delay10_q_net,
    q_12 => delay11_q_net,
    q_13 => delay12_q_net,
    q_14 => delay13_q_net,
    q_15 => delay14_q_net,
    q_16 => delay15_q_net
  );
  vector_slice : entity xil_defaultlib.psb3_0_vector_slice 
  port map (
    in_1 => mult0_p_net,
    in_2 => mult1_p_net,
    in_3 => mult2_p_net,
    in_4 => mult3_p_net,
    in_5 => mult4_p_net,
    in_6 => mult5_p_net,
    in_7 => mult6_p_net,
    in_8 => mult7_p_net,
    in_9 => mult8_p_net,
    in_10 => mult9_p_net,
    in_11 => mult10_p_net,
    in_12 => mult11_p_net,
    in_13 => mult12_p_net,
    in_14 => mult13_p_net,
    in_15 => mult14_p_net,
    in_16 => mult15_p_net,
    out_1 => slice0_y_net_x1,
    out_2 => slice1_y_net_x1,
    out_3 => slice2_y_net_x1,
    out_4 => slice3_y_net_x1,
    out_5 => slice4_y_net_x1,
    out_6 => slice5_y_net_x1,
    out_7 => slice6_y_net_x1,
    out_8 => slice7_y_net_x1,
    out_9 => slice8_y_net_x1,
    out_10 => slice9_y_net_x1,
    out_11 => slice10_y_net_x1,
    out_12 => slice11_y_net_x1,
    out_13 => slice12_y_net_x1,
    out_14 => slice13_y_net_x1,
    out_15 => slice14_y_net_x1,
    out_16 => slice15_y_net_x1
  );
  vector_slice1 : entity xil_defaultlib.psb3_0_vector_slice1 
  port map (
    in_1 => reinterpret0_output_port_net,
    in_2 => reinterpret1_output_port_net,
    in_3 => reinterpret2_output_port_net,
    in_4 => reinterpret3_output_port_net,
    in_5 => reinterpret4_output_port_net,
    in_6 => reinterpret5_output_port_net,
    in_7 => reinterpret6_output_port_net,
    in_8 => reinterpret7_output_port_net,
    in_9 => reinterpret8_output_port_net,
    in_10 => reinterpret9_output_port_net,
    in_11 => reinterpret10_output_port_net,
    in_12 => reinterpret11_output_port_net,
    in_13 => reinterpret12_output_port_net,
    in_14 => reinterpret13_output_port_net,
    in_15 => reinterpret14_output_port_net,
    in_16 => reinterpret15_output_port_net,
    out_1 => slice0_y_net_x0,
    out_2 => slice1_y_net_x0,
    out_3 => slice2_y_net_x0,
    out_4 => slice3_y_net_x0,
    out_5 => slice4_y_net_x0,
    out_6 => slice5_y_net_x0,
    out_7 => slice6_y_net_x0,
    out_8 => slice7_y_net_x0,
    out_9 => slice8_y_net_x0,
    out_10 => slice9_y_net_x0,
    out_11 => slice10_y_net_x0,
    out_12 => slice11_y_net_x0,
    out_13 => slice12_y_net_x0,
    out_14 => slice13_y_net_x0,
    out_15 => slice14_y_net_x0,
    out_16 => slice15_y_net_x0
  );
  vector_slice2 : entity xil_defaultlib.psb3_0_vector_slice2 
  port map (
    in_1 => addsub0_s_net,
    in_2 => addsub1_s_net,
    in_3 => addsub2_s_net,
    in_4 => addsub3_s_net,
    in_5 => addsub4_s_net,
    in_6 => addsub5_s_net,
    in_7 => addsub6_s_net,
    in_8 => addsub7_s_net,
    in_9 => addsub8_s_net,
    in_10 => addsub9_s_net,
    in_11 => addsub10_s_net,
    in_12 => addsub11_s_net,
    in_13 => addsub12_s_net,
    in_14 => addsub13_s_net,
    in_15 => addsub14_s_net,
    in_16 => addsub15_s_net,
    out_1 => slice0_y_net,
    out_2 => slice1_y_net,
    out_3 => slice2_y_net,
    out_4 => slice3_y_net,
    out_5 => slice4_y_net,
    out_6 => slice5_y_net,
    out_7 => slice6_y_net,
    out_8 => slice7_y_net,
    out_9 => slice8_y_net,
    out_10 => slice9_y_net,
    out_11 => slice10_y_net,
    out_12 => slice11_y_net,
    out_13 => slice12_y_net,
    out_14 => slice13_y_net,
    out_15 => slice14_y_net,
    out_16 => slice15_y_net
  );
  vector_to_scalar : entity xil_defaultlib.psb3_0_vector_to_scalar 
  port map (
    i_1 => delay0_q_net_x0,
    i_2 => delay1_q_net_x0,
    i_3 => delay2_q_net_x0,
    i_4 => delay3_q_net_x0,
    i_5 => delay4_q_net_x0,
    i_6 => delay5_q_net_x0,
    i_7 => delay6_q_net_x0,
    i_8 => delay7_q_net_x0,
    i_9 => delay8_q_net_x0,
    i_10 => delay9_q_net_x0,
    i_11 => delay10_q_net_x0,
    i_12 => delay11_q_net_x0,
    i_13 => delay12_q_net_x0,
    i_14 => delay13_q_net_x0,
    i_15 => delay14_q_net_x0,
    i_16 => delay15_q_net_x0,
    o => concat1_y_net_x1
  );
  vector_to_scalar1 : entity xil_defaultlib.psb3_0_vector_to_scalar1 
  port map (
    i_1 => delay0_q_net,
    i_2 => delay1_q_net,
    i_3 => delay2_q_net,
    i_4 => delay3_q_net,
    i_5 => delay4_q_net,
    i_6 => delay5_q_net,
    i_7 => delay6_q_net,
    i_8 => delay7_q_net,
    i_9 => delay8_q_net,
    i_10 => delay9_q_net,
    i_11 => delay10_q_net,
    i_12 => delay11_q_net,
    i_13 => delay12_q_net,
    i_14 => delay13_q_net,
    i_15 => delay14_q_net,
    i_16 => delay15_q_net,
    o => concat1_y_net_x0
  );
  vector_to_scalar2 : entity xil_defaultlib.psb3_0_vector_to_scalar2_x0 
  port map (
    i_1 => slice0_y_net,
    i_2 => slice1_y_net,
    i_3 => slice2_y_net,
    i_4 => slice3_y_net,
    i_5 => slice4_y_net,
    i_6 => slice5_y_net,
    i_7 => slice6_y_net,
    i_8 => slice7_y_net,
    i_9 => slice8_y_net,
    i_10 => slice9_y_net,
    i_11 => slice10_y_net,
    i_12 => slice11_y_net,
    i_13 => slice12_y_net,
    i_14 => slice13_y_net,
    i_15 => slice14_y_net,
    i_16 => slice15_y_net,
    o => concat1_y_net
  );
  constant17 : entity xil_defaultlib.sysgen_constant_71e89d757c 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant17_op_net
  );
  convert : entity xil_defaultlib.psb3_0_xlconvert 
  generic map (
    bool_conversion => 1,
    din_arith => 1,
    din_bin_pt => 0,
    din_width => 1,
    dout_arith => 1,
    dout_bin_pt => 0,
    dout_width => 1,
    latency => 1,
    overflow => xlWrap,
    quantization => xlTruncate
  )
  port map (
    clr => '0',
    en => "1",
    din => expression_dout_net,
    clk => clk_net,
    ce => ce_net,
    dout => convert_dout_net
  );
  expression : entity xil_defaultlib.sysgen_expr_7c83532765 
  port map (
    clr => '0',
    a => concat1_y_net_x1,
    b => concat1_y_net_x0,
    s => concat1_y_net,
    clk => clk_net,
    ce => ce_net,
    dout => expression_dout_net
  );
  register_x0 : entity xil_defaultlib.psb3_0_xlregister 
  generic map (
    d_width => 1,
    init_value => b"0"
  )
  port map (
    d => constant17_op_net,
    rst => gin_tl_reset_net,
    en => convert_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => register_q_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Overflow Detector add_im_2/Vector Delay
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_delay_x0 is
  port (
    d_1 : in std_logic_vector( 1-1 downto 0 );
    d_2 : in std_logic_vector( 1-1 downto 0 );
    d_3 : in std_logic_vector( 1-1 downto 0 );
    d_4 : in std_logic_vector( 1-1 downto 0 );
    d_5 : in std_logic_vector( 1-1 downto 0 );
    d_6 : in std_logic_vector( 1-1 downto 0 );
    d_7 : in std_logic_vector( 1-1 downto 0 );
    d_8 : in std_logic_vector( 1-1 downto 0 );
    d_9 : in std_logic_vector( 1-1 downto 0 );
    d_10 : in std_logic_vector( 1-1 downto 0 );
    d_11 : in std_logic_vector( 1-1 downto 0 );
    d_12 : in std_logic_vector( 1-1 downto 0 );
    d_13 : in std_logic_vector( 1-1 downto 0 );
    d_14 : in std_logic_vector( 1-1 downto 0 );
    d_15 : in std_logic_vector( 1-1 downto 0 );
    d_16 : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    q_1 : out std_logic_vector( 1-1 downto 0 );
    q_2 : out std_logic_vector( 1-1 downto 0 );
    q_3 : out std_logic_vector( 1-1 downto 0 );
    q_4 : out std_logic_vector( 1-1 downto 0 );
    q_5 : out std_logic_vector( 1-1 downto 0 );
    q_6 : out std_logic_vector( 1-1 downto 0 );
    q_7 : out std_logic_vector( 1-1 downto 0 );
    q_8 : out std_logic_vector( 1-1 downto 0 );
    q_9 : out std_logic_vector( 1-1 downto 0 );
    q_10 : out std_logic_vector( 1-1 downto 0 );
    q_11 : out std_logic_vector( 1-1 downto 0 );
    q_12 : out std_logic_vector( 1-1 downto 0 );
    q_13 : out std_logic_vector( 1-1 downto 0 );
    q_14 : out std_logic_vector( 1-1 downto 0 );
    q_15 : out std_logic_vector( 1-1 downto 0 );
    q_16 : out std_logic_vector( 1-1 downto 0 )
  );
end psb3_0_vector_delay_x0;
architecture structural of psb3_0_vector_delay_x0 is 
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay0_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay14_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay15_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay13_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay7_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay11_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay12_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay9_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay10_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal slice13_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal slice12_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 1-1 downto 0 );
begin
  q_1 <= delay0_q_net;
  q_2 <= delay1_q_net;
  q_3 <= delay2_q_net;
  q_4 <= delay3_q_net;
  q_5 <= delay4_q_net;
  q_6 <= delay5_q_net;
  q_7 <= delay6_q_net;
  q_8 <= delay7_q_net;
  q_9 <= delay8_q_net;
  q_10 <= delay9_q_net;
  q_11 <= delay10_q_net;
  q_12 <= delay11_q_net;
  q_13 <= delay12_q_net;
  q_14 <= delay13_q_net;
  q_15 <= delay14_q_net;
  q_16 <= delay15_q_net;
  slice0_y_net <= d_1;
  slice1_y_net <= d_2;
  slice2_y_net <= d_3;
  slice3_y_net <= d_4;
  slice4_y_net <= d_5;
  slice5_y_net <= d_6;
  slice6_y_net <= d_7;
  slice7_y_net <= d_8;
  slice8_y_net <= d_9;
  slice9_y_net <= d_10;
  slice10_y_net <= d_11;
  slice11_y_net <= d_12;
  slice12_y_net <= d_13;
  slice13_y_net <= d_14;
  slice14_y_net <= d_15;
  slice15_y_net <= d_16;
  clk_net <= clk_1;
  ce_net <= ce_1;
  delay0 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice0_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay0_q_net
  );
  delay1 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice2_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay3 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice3_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  delay4 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice4_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net
  );
  delay5 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice5_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  delay6 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice6_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay6_q_net
  );
  delay7 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice7_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay7_q_net
  );
  delay8 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice8_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay8_q_net
  );
  delay9 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice9_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay9_q_net
  );
  delay10 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice10_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay10_q_net
  );
  delay11 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice11_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay11_q_net
  );
  delay12 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice12_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay12_q_net
  );
  delay13 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice13_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay13_q_net
  );
  delay14 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice14_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay14_q_net
  );
  delay15 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice15_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay15_q_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Overflow Detector add_im_2/Vector Delay1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_delay1_x0 is
  port (
    d_1 : in std_logic_vector( 1-1 downto 0 );
    d_2 : in std_logic_vector( 1-1 downto 0 );
    d_3 : in std_logic_vector( 1-1 downto 0 );
    d_4 : in std_logic_vector( 1-1 downto 0 );
    d_5 : in std_logic_vector( 1-1 downto 0 );
    d_6 : in std_logic_vector( 1-1 downto 0 );
    d_7 : in std_logic_vector( 1-1 downto 0 );
    d_8 : in std_logic_vector( 1-1 downto 0 );
    d_9 : in std_logic_vector( 1-1 downto 0 );
    d_10 : in std_logic_vector( 1-1 downto 0 );
    d_11 : in std_logic_vector( 1-1 downto 0 );
    d_12 : in std_logic_vector( 1-1 downto 0 );
    d_13 : in std_logic_vector( 1-1 downto 0 );
    d_14 : in std_logic_vector( 1-1 downto 0 );
    d_15 : in std_logic_vector( 1-1 downto 0 );
    d_16 : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    q_1 : out std_logic_vector( 1-1 downto 0 );
    q_2 : out std_logic_vector( 1-1 downto 0 );
    q_3 : out std_logic_vector( 1-1 downto 0 );
    q_4 : out std_logic_vector( 1-1 downto 0 );
    q_5 : out std_logic_vector( 1-1 downto 0 );
    q_6 : out std_logic_vector( 1-1 downto 0 );
    q_7 : out std_logic_vector( 1-1 downto 0 );
    q_8 : out std_logic_vector( 1-1 downto 0 );
    q_9 : out std_logic_vector( 1-1 downto 0 );
    q_10 : out std_logic_vector( 1-1 downto 0 );
    q_11 : out std_logic_vector( 1-1 downto 0 );
    q_12 : out std_logic_vector( 1-1 downto 0 );
    q_13 : out std_logic_vector( 1-1 downto 0 );
    q_14 : out std_logic_vector( 1-1 downto 0 );
    q_15 : out std_logic_vector( 1-1 downto 0 );
    q_16 : out std_logic_vector( 1-1 downto 0 )
  );
end psb3_0_vector_delay1_x0;
architecture structural of psb3_0_vector_delay1_x0 is 
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay0_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay9_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay15_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay12_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay13_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay10_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay7_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal slice9_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay14_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal slice0_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay11_q_net : std_logic_vector( 1-1 downto 0 );
begin
  q_1 <= delay0_q_net;
  q_2 <= delay1_q_net;
  q_3 <= delay2_q_net;
  q_4 <= delay3_q_net;
  q_5 <= delay4_q_net;
  q_6 <= delay5_q_net;
  q_7 <= delay6_q_net;
  q_8 <= delay7_q_net;
  q_9 <= delay8_q_net;
  q_10 <= delay9_q_net;
  q_11 <= delay10_q_net;
  q_12 <= delay11_q_net;
  q_13 <= delay12_q_net;
  q_14 <= delay13_q_net;
  q_15 <= delay14_q_net;
  q_16 <= delay15_q_net;
  slice0_y_net <= d_1;
  slice1_y_net <= d_2;
  slice2_y_net <= d_3;
  slice3_y_net <= d_4;
  slice4_y_net <= d_5;
  slice5_y_net <= d_6;
  slice6_y_net <= d_7;
  slice7_y_net <= d_8;
  slice8_y_net <= d_9;
  slice9_y_net <= d_10;
  slice10_y_net <= d_11;
  slice11_y_net <= d_12;
  slice12_y_net <= d_13;
  slice13_y_net <= d_14;
  slice14_y_net <= d_15;
  slice15_y_net <= d_16;
  clk_net <= clk_1;
  ce_net <= ce_1;
  delay0 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice0_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay0_q_net
  );
  delay1 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice2_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay3 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice3_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  delay4 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice4_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net
  );
  delay5 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice5_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  delay6 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice6_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay6_q_net
  );
  delay7 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice7_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay7_q_net
  );
  delay8 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice8_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay8_q_net
  );
  delay9 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice9_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay9_q_net
  );
  delay10 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice10_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay10_q_net
  );
  delay11 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice11_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay11_q_net
  );
  delay12 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice12_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay12_q_net
  );
  delay13 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice13_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay13_q_net
  );
  delay14 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice14_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay14_q_net
  );
  delay15 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice15_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay15_q_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Overflow Detector add_im_2/Vector Slice
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_slice_x0 is
  port (
    in_1 : in std_logic_vector( 16-1 downto 0 );
    in_2 : in std_logic_vector( 16-1 downto 0 );
    in_3 : in std_logic_vector( 16-1 downto 0 );
    in_4 : in std_logic_vector( 16-1 downto 0 );
    in_5 : in std_logic_vector( 16-1 downto 0 );
    in_6 : in std_logic_vector( 16-1 downto 0 );
    in_7 : in std_logic_vector( 16-1 downto 0 );
    in_8 : in std_logic_vector( 16-1 downto 0 );
    in_9 : in std_logic_vector( 16-1 downto 0 );
    in_10 : in std_logic_vector( 16-1 downto 0 );
    in_11 : in std_logic_vector( 16-1 downto 0 );
    in_12 : in std_logic_vector( 16-1 downto 0 );
    in_13 : in std_logic_vector( 16-1 downto 0 );
    in_14 : in std_logic_vector( 16-1 downto 0 );
    in_15 : in std_logic_vector( 16-1 downto 0 );
    in_16 : in std_logic_vector( 16-1 downto 0 );
    out_1 : out std_logic_vector( 1-1 downto 0 );
    out_2 : out std_logic_vector( 1-1 downto 0 );
    out_3 : out std_logic_vector( 1-1 downto 0 );
    out_4 : out std_logic_vector( 1-1 downto 0 );
    out_5 : out std_logic_vector( 1-1 downto 0 );
    out_6 : out std_logic_vector( 1-1 downto 0 );
    out_7 : out std_logic_vector( 1-1 downto 0 );
    out_8 : out std_logic_vector( 1-1 downto 0 );
    out_9 : out std_logic_vector( 1-1 downto 0 );
    out_10 : out std_logic_vector( 1-1 downto 0 );
    out_11 : out std_logic_vector( 1-1 downto 0 );
    out_12 : out std_logic_vector( 1-1 downto 0 );
    out_13 : out std_logic_vector( 1-1 downto 0 );
    out_14 : out std_logic_vector( 1-1 downto 0 );
    out_15 : out std_logic_vector( 1-1 downto 0 );
    out_16 : out std_logic_vector( 1-1 downto 0 )
  );
end psb3_0_vector_slice_x0;
architecture structural of psb3_0_vector_slice_x0 is 
  signal slice9_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 1-1 downto 0 );
  signal mult0_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult1_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult2_p_net : std_logic_vector( 16-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 1-1 downto 0 );
  signal mult3_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult8_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult7_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult13_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult12_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult6_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult5_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult15_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult4_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult9_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult10_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult14_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult11_p_net : std_logic_vector( 16-1 downto 0 );
begin
  out_1 <= slice0_y_net;
  out_2 <= slice1_y_net;
  out_3 <= slice2_y_net;
  out_4 <= slice3_y_net;
  out_5 <= slice4_y_net;
  out_6 <= slice5_y_net;
  out_7 <= slice6_y_net;
  out_8 <= slice7_y_net;
  out_9 <= slice8_y_net;
  out_10 <= slice9_y_net;
  out_11 <= slice10_y_net;
  out_12 <= slice11_y_net;
  out_13 <= slice12_y_net;
  out_14 <= slice13_y_net;
  out_15 <= slice14_y_net;
  out_16 <= slice15_y_net;
  mult0_p_net <= in_1;
  mult1_p_net <= in_2;
  mult2_p_net <= in_3;
  mult3_p_net <= in_4;
  mult4_p_net <= in_5;
  mult5_p_net <= in_6;
  mult6_p_net <= in_7;
  mult7_p_net <= in_8;
  mult8_p_net <= in_9;
  mult9_p_net <= in_10;
  mult10_p_net <= in_11;
  mult11_p_net <= in_12;
  mult12_p_net <= in_13;
  mult13_p_net <= in_14;
  mult14_p_net <= in_15;
  mult15_p_net <= in_16;
  slice0 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult0_p_net,
    y => slice0_y_net
  );
  slice1 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult1_p_net,
    y => slice1_y_net
  );
  slice2 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult2_p_net,
    y => slice2_y_net
  );
  slice3 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult3_p_net,
    y => slice3_y_net
  );
  slice4 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult4_p_net,
    y => slice4_y_net
  );
  slice5 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult5_p_net,
    y => slice5_y_net
  );
  slice6 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult6_p_net,
    y => slice6_y_net
  );
  slice7 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult7_p_net,
    y => slice7_y_net
  );
  slice8 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult8_p_net,
    y => slice8_y_net
  );
  slice9 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult9_p_net,
    y => slice9_y_net
  );
  slice10 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult10_p_net,
    y => slice10_y_net
  );
  slice11 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult11_p_net,
    y => slice11_y_net
  );
  slice12 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult12_p_net,
    y => slice12_y_net
  );
  slice13 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult13_p_net,
    y => slice13_y_net
  );
  slice14 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult14_p_net,
    y => slice14_y_net
  );
  slice15 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult15_p_net,
    y => slice15_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Overflow Detector add_im_2/Vector Slice1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_slice1_x0 is
  port (
    in_1 : in std_logic_vector( 16-1 downto 0 );
    in_2 : in std_logic_vector( 16-1 downto 0 );
    in_3 : in std_logic_vector( 16-1 downto 0 );
    in_4 : in std_logic_vector( 16-1 downto 0 );
    in_5 : in std_logic_vector( 16-1 downto 0 );
    in_6 : in std_logic_vector( 16-1 downto 0 );
    in_7 : in std_logic_vector( 16-1 downto 0 );
    in_8 : in std_logic_vector( 16-1 downto 0 );
    in_9 : in std_logic_vector( 16-1 downto 0 );
    in_10 : in std_logic_vector( 16-1 downto 0 );
    in_11 : in std_logic_vector( 16-1 downto 0 );
    in_12 : in std_logic_vector( 16-1 downto 0 );
    in_13 : in std_logic_vector( 16-1 downto 0 );
    in_14 : in std_logic_vector( 16-1 downto 0 );
    in_15 : in std_logic_vector( 16-1 downto 0 );
    in_16 : in std_logic_vector( 16-1 downto 0 );
    out_1 : out std_logic_vector( 1-1 downto 0 );
    out_2 : out std_logic_vector( 1-1 downto 0 );
    out_3 : out std_logic_vector( 1-1 downto 0 );
    out_4 : out std_logic_vector( 1-1 downto 0 );
    out_5 : out std_logic_vector( 1-1 downto 0 );
    out_6 : out std_logic_vector( 1-1 downto 0 );
    out_7 : out std_logic_vector( 1-1 downto 0 );
    out_8 : out std_logic_vector( 1-1 downto 0 );
    out_9 : out std_logic_vector( 1-1 downto 0 );
    out_10 : out std_logic_vector( 1-1 downto 0 );
    out_11 : out std_logic_vector( 1-1 downto 0 );
    out_12 : out std_logic_vector( 1-1 downto 0 );
    out_13 : out std_logic_vector( 1-1 downto 0 );
    out_14 : out std_logic_vector( 1-1 downto 0 );
    out_15 : out std_logic_vector( 1-1 downto 0 );
    out_16 : out std_logic_vector( 1-1 downto 0 )
  );
end psb3_0_vector_slice1_x0;
architecture structural of psb3_0_vector_slice1_x0 is 
  signal slice1_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
begin
  out_1 <= slice0_y_net;
  out_2 <= slice1_y_net;
  out_3 <= slice2_y_net;
  out_4 <= slice3_y_net;
  out_5 <= slice4_y_net;
  out_6 <= slice5_y_net;
  out_7 <= slice6_y_net;
  out_8 <= slice7_y_net;
  out_9 <= slice8_y_net;
  out_10 <= slice9_y_net;
  out_11 <= slice10_y_net;
  out_12 <= slice11_y_net;
  out_13 <= slice12_y_net;
  out_14 <= slice13_y_net;
  out_15 <= slice14_y_net;
  out_16 <= slice15_y_net;
  reinterpret0_output_port_net <= in_1;
  reinterpret1_output_port_net <= in_2;
  reinterpret2_output_port_net <= in_3;
  reinterpret3_output_port_net <= in_4;
  reinterpret4_output_port_net <= in_5;
  reinterpret5_output_port_net <= in_6;
  reinterpret6_output_port_net <= in_7;
  reinterpret7_output_port_net <= in_8;
  reinterpret8_output_port_net <= in_9;
  reinterpret9_output_port_net <= in_10;
  reinterpret10_output_port_net <= in_11;
  reinterpret11_output_port_net <= in_12;
  reinterpret12_output_port_net <= in_13;
  reinterpret13_output_port_net <= in_14;
  reinterpret14_output_port_net <= in_15;
  reinterpret15_output_port_net <= in_16;
  slice0 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret0_output_port_net,
    y => slice0_y_net
  );
  slice1 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret1_output_port_net,
    y => slice1_y_net
  );
  slice2 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret2_output_port_net,
    y => slice2_y_net
  );
  slice3 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret3_output_port_net,
    y => slice3_y_net
  );
  slice4 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret4_output_port_net,
    y => slice4_y_net
  );
  slice5 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret5_output_port_net,
    y => slice5_y_net
  );
  slice6 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret6_output_port_net,
    y => slice6_y_net
  );
  slice7 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret7_output_port_net,
    y => slice7_y_net
  );
  slice8 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret8_output_port_net,
    y => slice8_y_net
  );
  slice9 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret9_output_port_net,
    y => slice9_y_net
  );
  slice10 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret10_output_port_net,
    y => slice10_y_net
  );
  slice11 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret11_output_port_net,
    y => slice11_y_net
  );
  slice12 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret12_output_port_net,
    y => slice12_y_net
  );
  slice13 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret13_output_port_net,
    y => slice13_y_net
  );
  slice14 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret14_output_port_net,
    y => slice14_y_net
  );
  slice15 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret15_output_port_net,
    y => slice15_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Overflow Detector add_im_2/Vector Slice2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_slice2_x0 is
  port (
    in_1 : in std_logic_vector( 16-1 downto 0 );
    in_2 : in std_logic_vector( 16-1 downto 0 );
    in_3 : in std_logic_vector( 16-1 downto 0 );
    in_4 : in std_logic_vector( 16-1 downto 0 );
    in_5 : in std_logic_vector( 16-1 downto 0 );
    in_6 : in std_logic_vector( 16-1 downto 0 );
    in_7 : in std_logic_vector( 16-1 downto 0 );
    in_8 : in std_logic_vector( 16-1 downto 0 );
    in_9 : in std_logic_vector( 16-1 downto 0 );
    in_10 : in std_logic_vector( 16-1 downto 0 );
    in_11 : in std_logic_vector( 16-1 downto 0 );
    in_12 : in std_logic_vector( 16-1 downto 0 );
    in_13 : in std_logic_vector( 16-1 downto 0 );
    in_14 : in std_logic_vector( 16-1 downto 0 );
    in_15 : in std_logic_vector( 16-1 downto 0 );
    in_16 : in std_logic_vector( 16-1 downto 0 );
    out_1 : out std_logic_vector( 1-1 downto 0 );
    out_2 : out std_logic_vector( 1-1 downto 0 );
    out_3 : out std_logic_vector( 1-1 downto 0 );
    out_4 : out std_logic_vector( 1-1 downto 0 );
    out_5 : out std_logic_vector( 1-1 downto 0 );
    out_6 : out std_logic_vector( 1-1 downto 0 );
    out_7 : out std_logic_vector( 1-1 downto 0 );
    out_8 : out std_logic_vector( 1-1 downto 0 );
    out_9 : out std_logic_vector( 1-1 downto 0 );
    out_10 : out std_logic_vector( 1-1 downto 0 );
    out_11 : out std_logic_vector( 1-1 downto 0 );
    out_12 : out std_logic_vector( 1-1 downto 0 );
    out_13 : out std_logic_vector( 1-1 downto 0 );
    out_14 : out std_logic_vector( 1-1 downto 0 );
    out_15 : out std_logic_vector( 1-1 downto 0 );
    out_16 : out std_logic_vector( 1-1 downto 0 )
  );
end psb3_0_vector_slice2_x0;
architecture structural of psb3_0_vector_slice2_x0 is 
  signal addsub0_s_net : std_logic_vector( 16-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 1-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub6_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub5_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub8_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub13_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub12_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub3_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub9_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub7_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub10_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub14_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub11_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub15_s_net : std_logic_vector( 16-1 downto 0 );
begin
  out_1 <= slice0_y_net;
  out_2 <= slice1_y_net;
  out_3 <= slice2_y_net;
  out_4 <= slice3_y_net;
  out_5 <= slice4_y_net;
  out_6 <= slice5_y_net;
  out_7 <= slice6_y_net;
  out_8 <= slice7_y_net;
  out_9 <= slice8_y_net;
  out_10 <= slice9_y_net;
  out_11 <= slice10_y_net;
  out_12 <= slice11_y_net;
  out_13 <= slice12_y_net;
  out_14 <= slice13_y_net;
  out_15 <= slice14_y_net;
  out_16 <= slice15_y_net;
  addsub0_s_net <= in_1;
  addsub1_s_net <= in_2;
  addsub2_s_net <= in_3;
  addsub3_s_net <= in_4;
  addsub4_s_net <= in_5;
  addsub5_s_net <= in_6;
  addsub6_s_net <= in_7;
  addsub7_s_net <= in_8;
  addsub8_s_net <= in_9;
  addsub9_s_net <= in_10;
  addsub10_s_net <= in_11;
  addsub11_s_net <= in_12;
  addsub12_s_net <= in_13;
  addsub13_s_net <= in_14;
  addsub14_s_net <= in_15;
  addsub15_s_net <= in_16;
  slice0 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub0_s_net,
    y => slice0_y_net
  );
  slice1 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub1_s_net,
    y => slice1_y_net
  );
  slice2 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub2_s_net,
    y => slice2_y_net
  );
  slice3 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub3_s_net,
    y => slice3_y_net
  );
  slice4 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub4_s_net,
    y => slice4_y_net
  );
  slice5 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub5_s_net,
    y => slice5_y_net
  );
  slice6 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub6_s_net,
    y => slice6_y_net
  );
  slice7 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub7_s_net,
    y => slice7_y_net
  );
  slice8 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub8_s_net,
    y => slice8_y_net
  );
  slice9 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub9_s_net,
    y => slice9_y_net
  );
  slice10 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub10_s_net,
    y => slice10_y_net
  );
  slice11 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub11_s_net,
    y => slice11_y_net
  );
  slice12 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub12_s_net,
    y => slice12_y_net
  );
  slice13 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub13_s_net,
    y => slice13_y_net
  );
  slice14 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub14_s_net,
    y => slice14_y_net
  );
  slice15 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub15_s_net,
    y => slice15_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Overflow Detector add_im_2/Vector to Scalar
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_to_scalar_x0 is
  port (
    i_1 : in std_logic_vector( 1-1 downto 0 );
    i_2 : in std_logic_vector( 1-1 downto 0 );
    i_3 : in std_logic_vector( 1-1 downto 0 );
    i_4 : in std_logic_vector( 1-1 downto 0 );
    i_5 : in std_logic_vector( 1-1 downto 0 );
    i_6 : in std_logic_vector( 1-1 downto 0 );
    i_7 : in std_logic_vector( 1-1 downto 0 );
    i_8 : in std_logic_vector( 1-1 downto 0 );
    i_9 : in std_logic_vector( 1-1 downto 0 );
    i_10 : in std_logic_vector( 1-1 downto 0 );
    i_11 : in std_logic_vector( 1-1 downto 0 );
    i_12 : in std_logic_vector( 1-1 downto 0 );
    i_13 : in std_logic_vector( 1-1 downto 0 );
    i_14 : in std_logic_vector( 1-1 downto 0 );
    i_15 : in std_logic_vector( 1-1 downto 0 );
    i_16 : in std_logic_vector( 1-1 downto 0 );
    o : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_vector_to_scalar_x0;
architecture structural of psb3_0_vector_to_scalar_x0 is 
  signal concat1_y_net : std_logic_vector( 16-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay7_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay15_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay11_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay10_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay12_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay14_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay0_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay9_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay13_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
begin
  o <= concat1_y_net;
  delay0_q_net <= i_1;
  delay1_q_net <= i_2;
  delay2_q_net <= i_3;
  delay3_q_net <= i_4;
  delay4_q_net <= i_5;
  delay5_q_net <= i_6;
  delay6_q_net <= i_7;
  delay7_q_net <= i_8;
  delay8_q_net <= i_9;
  delay9_q_net <= i_10;
  delay10_q_net <= i_11;
  delay11_q_net <= i_12;
  delay12_q_net <= i_13;
  delay13_q_net <= i_14;
  delay14_q_net <= i_15;
  delay15_q_net <= i_16;
  concat1 : entity xil_defaultlib.sysgen_concat_d977c66e35 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => delay15_q_net,
    in1 => delay14_q_net,
    in2 => delay13_q_net,
    in3 => delay12_q_net,
    in4 => delay11_q_net,
    in5 => delay10_q_net,
    in6 => delay9_q_net,
    in7 => delay8_q_net,
    in8 => delay7_q_net,
    in9 => delay6_q_net,
    in10 => delay5_q_net,
    in11 => delay4_q_net,
    in12 => delay3_q_net,
    in13 => delay2_q_net,
    in14 => delay1_q_net,
    in15 => delay0_q_net,
    y => concat1_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Overflow Detector add_im_2/Vector to Scalar1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_to_scalar1_x0 is
  port (
    i_1 : in std_logic_vector( 1-1 downto 0 );
    i_2 : in std_logic_vector( 1-1 downto 0 );
    i_3 : in std_logic_vector( 1-1 downto 0 );
    i_4 : in std_logic_vector( 1-1 downto 0 );
    i_5 : in std_logic_vector( 1-1 downto 0 );
    i_6 : in std_logic_vector( 1-1 downto 0 );
    i_7 : in std_logic_vector( 1-1 downto 0 );
    i_8 : in std_logic_vector( 1-1 downto 0 );
    i_9 : in std_logic_vector( 1-1 downto 0 );
    i_10 : in std_logic_vector( 1-1 downto 0 );
    i_11 : in std_logic_vector( 1-1 downto 0 );
    i_12 : in std_logic_vector( 1-1 downto 0 );
    i_13 : in std_logic_vector( 1-1 downto 0 );
    i_14 : in std_logic_vector( 1-1 downto 0 );
    i_15 : in std_logic_vector( 1-1 downto 0 );
    i_16 : in std_logic_vector( 1-1 downto 0 );
    o : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_vector_to_scalar1_x0;
architecture structural of psb3_0_vector_to_scalar1_x0 is 
  signal concat1_y_net : std_logic_vector( 16-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay0_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay10_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay11_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay9_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay13_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay12_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay14_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay15_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay7_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 1-1 downto 0 );
begin
  o <= concat1_y_net;
  delay0_q_net <= i_1;
  delay1_q_net <= i_2;
  delay2_q_net <= i_3;
  delay3_q_net <= i_4;
  delay4_q_net <= i_5;
  delay5_q_net <= i_6;
  delay6_q_net <= i_7;
  delay7_q_net <= i_8;
  delay8_q_net <= i_9;
  delay9_q_net <= i_10;
  delay10_q_net <= i_11;
  delay11_q_net <= i_12;
  delay12_q_net <= i_13;
  delay13_q_net <= i_14;
  delay14_q_net <= i_15;
  delay15_q_net <= i_16;
  concat1 : entity xil_defaultlib.sysgen_concat_d977c66e35 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => delay15_q_net,
    in1 => delay14_q_net,
    in2 => delay13_q_net,
    in3 => delay12_q_net,
    in4 => delay11_q_net,
    in5 => delay10_q_net,
    in6 => delay9_q_net,
    in7 => delay8_q_net,
    in8 => delay7_q_net,
    in9 => delay6_q_net,
    in10 => delay5_q_net,
    in11 => delay4_q_net,
    in12 => delay3_q_net,
    in13 => delay2_q_net,
    in14 => delay1_q_net,
    in15 => delay0_q_net,
    y => concat1_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Overflow Detector add_im_2/Vector to Scalar2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_to_scalar2_x1 is
  port (
    i_1 : in std_logic_vector( 1-1 downto 0 );
    i_2 : in std_logic_vector( 1-1 downto 0 );
    i_3 : in std_logic_vector( 1-1 downto 0 );
    i_4 : in std_logic_vector( 1-1 downto 0 );
    i_5 : in std_logic_vector( 1-1 downto 0 );
    i_6 : in std_logic_vector( 1-1 downto 0 );
    i_7 : in std_logic_vector( 1-1 downto 0 );
    i_8 : in std_logic_vector( 1-1 downto 0 );
    i_9 : in std_logic_vector( 1-1 downto 0 );
    i_10 : in std_logic_vector( 1-1 downto 0 );
    i_11 : in std_logic_vector( 1-1 downto 0 );
    i_12 : in std_logic_vector( 1-1 downto 0 );
    i_13 : in std_logic_vector( 1-1 downto 0 );
    i_14 : in std_logic_vector( 1-1 downto 0 );
    i_15 : in std_logic_vector( 1-1 downto 0 );
    i_16 : in std_logic_vector( 1-1 downto 0 );
    o : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_vector_to_scalar2_x1;
architecture structural of psb3_0_vector_to_scalar2_x1 is 
  signal concat1_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 1-1 downto 0 );
begin
  o <= concat1_y_net;
  slice0_y_net <= i_1;
  slice1_y_net <= i_2;
  slice2_y_net <= i_3;
  slice3_y_net <= i_4;
  slice4_y_net <= i_5;
  slice5_y_net <= i_6;
  slice6_y_net <= i_7;
  slice7_y_net <= i_8;
  slice8_y_net <= i_9;
  slice9_y_net <= i_10;
  slice10_y_net <= i_11;
  slice11_y_net <= i_12;
  slice12_y_net <= i_13;
  slice13_y_net <= i_14;
  slice14_y_net <= i_15;
  slice15_y_net <= i_16;
  concat1 : entity xil_defaultlib.sysgen_concat_d977c66e35 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => slice15_y_net,
    in1 => slice14_y_net,
    in2 => slice13_y_net,
    in3 => slice12_y_net,
    in4 => slice11_y_net,
    in5 => slice10_y_net,
    in6 => slice9_y_net,
    in7 => slice8_y_net,
    in8 => slice7_y_net,
    in9 => slice6_y_net,
    in10 => slice5_y_net,
    in11 => slice4_y_net,
    in12 => slice3_y_net,
    in13 => slice2_y_net,
    in14 => slice1_y_net,
    in15 => slice0_y_net,
    y => concat1_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Overflow Detector add_im_2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_overflow_detector_add_im_2 is
  port (
    rst : in std_logic_vector( 1-1 downto 0 );
    a_1 : in std_logic_vector( 16-1 downto 0 );
    b_1 : in std_logic_vector( 16-1 downto 0 );
    s_1 : in std_logic_vector( 16-1 downto 0 );
    a_2 : in std_logic_vector( 16-1 downto 0 );
    a_3 : in std_logic_vector( 16-1 downto 0 );
    a_4 : in std_logic_vector( 16-1 downto 0 );
    a_5 : in std_logic_vector( 16-1 downto 0 );
    a_6 : in std_logic_vector( 16-1 downto 0 );
    a_7 : in std_logic_vector( 16-1 downto 0 );
    a_8 : in std_logic_vector( 16-1 downto 0 );
    a_9 : in std_logic_vector( 16-1 downto 0 );
    a_10 : in std_logic_vector( 16-1 downto 0 );
    a_11 : in std_logic_vector( 16-1 downto 0 );
    a_12 : in std_logic_vector( 16-1 downto 0 );
    a_13 : in std_logic_vector( 16-1 downto 0 );
    a_14 : in std_logic_vector( 16-1 downto 0 );
    a_15 : in std_logic_vector( 16-1 downto 0 );
    a_16 : in std_logic_vector( 16-1 downto 0 );
    b_2 : in std_logic_vector( 16-1 downto 0 );
    b_3 : in std_logic_vector( 16-1 downto 0 );
    b_4 : in std_logic_vector( 16-1 downto 0 );
    b_5 : in std_logic_vector( 16-1 downto 0 );
    b_6 : in std_logic_vector( 16-1 downto 0 );
    b_7 : in std_logic_vector( 16-1 downto 0 );
    b_8 : in std_logic_vector( 16-1 downto 0 );
    b_9 : in std_logic_vector( 16-1 downto 0 );
    b_10 : in std_logic_vector( 16-1 downto 0 );
    b_11 : in std_logic_vector( 16-1 downto 0 );
    b_12 : in std_logic_vector( 16-1 downto 0 );
    b_13 : in std_logic_vector( 16-1 downto 0 );
    b_14 : in std_logic_vector( 16-1 downto 0 );
    b_15 : in std_logic_vector( 16-1 downto 0 );
    b_16 : in std_logic_vector( 16-1 downto 0 );
    s_2 : in std_logic_vector( 16-1 downto 0 );
    s_3 : in std_logic_vector( 16-1 downto 0 );
    s_4 : in std_logic_vector( 16-1 downto 0 );
    s_5 : in std_logic_vector( 16-1 downto 0 );
    s_6 : in std_logic_vector( 16-1 downto 0 );
    s_7 : in std_logic_vector( 16-1 downto 0 );
    s_8 : in std_logic_vector( 16-1 downto 0 );
    s_9 : in std_logic_vector( 16-1 downto 0 );
    s_10 : in std_logic_vector( 16-1 downto 0 );
    s_11 : in std_logic_vector( 16-1 downto 0 );
    s_12 : in std_logic_vector( 16-1 downto 0 );
    s_13 : in std_logic_vector( 16-1 downto 0 );
    s_14 : in std_logic_vector( 16-1 downto 0 );
    s_15 : in std_logic_vector( 16-1 downto 0 );
    s_16 : in std_logic_vector( 16-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    ov : out std_logic_vector( 1-1 downto 0 )
  );
end psb3_0_overflow_detector_add_im_2;
architecture structural of psb3_0_overflow_detector_add_im_2 is 
  signal mult4_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult5_p_net : std_logic_vector( 16-1 downto 0 );
  signal addsub0_s_net : std_logic_vector( 16-1 downto 0 );
  signal mult2_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult0_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult1_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult3_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult7_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult6_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult8_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult9_p_net : std_logic_vector( 16-1 downto 0 );
  signal register_q_net : std_logic_vector( 1-1 downto 0 );
  signal gin_tl_reset_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub3_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub5_s_net : std_logic_vector( 16-1 downto 0 );
  signal mult12_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub6_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub8_s_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub9_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub11_s_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mult15_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mult10_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub7_s_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub10_s_net : std_logic_vector( 16-1 downto 0 );
  signal mult13_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult11_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 16-1 downto 0 );
  signal mult14_p_net : std_logic_vector( 16-1 downto 0 );
  signal delay2_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay5_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay13_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice3_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal slice7_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice9_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal slice5_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal delay13_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay14_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice10_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal slice12_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal slice13_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay7_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice14_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal delay15_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice0_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice2_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay0_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay8_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay4_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay11_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay14_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay7_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal addsub15_s_net : std_logic_vector( 16-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal delay10_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay12_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice1_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice3_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay15_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice4_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal delay3_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal addsub14_s_net : std_logic_vector( 16-1 downto 0 );
  signal delay6_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay9_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice0_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal slice6_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal slice11_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal slice2_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal delay10_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice1_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal delay0_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay12_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice4_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal slice8_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal slice15_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal addsub12_s_net : std_logic_vector( 16-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay9_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay11_q_net : std_logic_vector( 1-1 downto 0 );
  signal addsub13_s_net : std_logic_vector( 16-1 downto 0 );
  signal concat1_y_net_x1 : std_logic_vector( 16-1 downto 0 );
  signal slice12_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice11_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice7_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice13_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice14_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice9_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 1-1 downto 0 );
  signal concat1_y_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal slice6_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice8_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice15_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 1-1 downto 0 );
  signal constant17_op_net : std_logic_vector( 1-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 1-1 downto 0 );
  signal concat1_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 1-1 downto 0 );
  signal convert_dout_net : std_logic_vector( 1-1 downto 0 );
  signal expression_dout_net : std_logic_vector( 1-1 downto 0 );
  signal slice5_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice10_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 1-1 downto 0 );
begin
  ov <= register_q_net;
  gin_tl_reset_net <= rst;
  mult0_p_net <= a_1;
  reinterpret0_output_port_net <= b_1;
  addsub0_s_net <= s_1;
  mult1_p_net <= a_2;
  mult2_p_net <= a_3;
  mult3_p_net <= a_4;
  mult4_p_net <= a_5;
  mult5_p_net <= a_6;
  mult6_p_net <= a_7;
  mult7_p_net <= a_8;
  mult8_p_net <= a_9;
  mult9_p_net <= a_10;
  mult10_p_net <= a_11;
  mult11_p_net <= a_12;
  mult12_p_net <= a_13;
  mult13_p_net <= a_14;
  mult14_p_net <= a_15;
  mult15_p_net <= a_16;
  reinterpret1_output_port_net <= b_2;
  reinterpret2_output_port_net <= b_3;
  reinterpret3_output_port_net <= b_4;
  reinterpret4_output_port_net <= b_5;
  reinterpret5_output_port_net <= b_6;
  reinterpret6_output_port_net <= b_7;
  reinterpret7_output_port_net <= b_8;
  reinterpret8_output_port_net <= b_9;
  reinterpret9_output_port_net <= b_10;
  reinterpret10_output_port_net <= b_11;
  reinterpret11_output_port_net <= b_12;
  reinterpret12_output_port_net <= b_13;
  reinterpret13_output_port_net <= b_14;
  reinterpret14_output_port_net <= b_15;
  reinterpret15_output_port_net <= b_16;
  addsub1_s_net <= s_2;
  addsub2_s_net <= s_3;
  addsub3_s_net <= s_4;
  addsub4_s_net <= s_5;
  addsub5_s_net <= s_6;
  addsub6_s_net <= s_7;
  addsub7_s_net <= s_8;
  addsub8_s_net <= s_9;
  addsub9_s_net <= s_10;
  addsub10_s_net <= s_11;
  addsub11_s_net <= s_12;
  addsub12_s_net <= s_13;
  addsub13_s_net <= s_14;
  addsub14_s_net <= s_15;
  addsub15_s_net <= s_16;
  clk_net <= clk_1;
  ce_net <= ce_1;
  vector_delay : entity xil_defaultlib.psb3_0_vector_delay_x0 
  port map (
    d_1 => slice0_y_net_x1,
    d_2 => slice1_y_net_x1,
    d_3 => slice2_y_net_x1,
    d_4 => slice3_y_net_x1,
    d_5 => slice4_y_net_x1,
    d_6 => slice5_y_net_x1,
    d_7 => slice6_y_net_x1,
    d_8 => slice7_y_net_x1,
    d_9 => slice8_y_net_x1,
    d_10 => slice9_y_net_x1,
    d_11 => slice10_y_net_x1,
    d_12 => slice11_y_net_x1,
    d_13 => slice12_y_net_x1,
    d_14 => slice13_y_net_x1,
    d_15 => slice14_y_net_x1,
    d_16 => slice15_y_net_x1,
    clk_1 => clk_net,
    ce_1 => ce_net,
    q_1 => delay0_q_net_x0,
    q_2 => delay1_q_net_x0,
    q_3 => delay2_q_net_x0,
    q_4 => delay3_q_net_x0,
    q_5 => delay4_q_net_x0,
    q_6 => delay5_q_net_x0,
    q_7 => delay6_q_net_x0,
    q_8 => delay7_q_net_x0,
    q_9 => delay8_q_net_x0,
    q_10 => delay9_q_net_x0,
    q_11 => delay10_q_net_x0,
    q_12 => delay11_q_net_x0,
    q_13 => delay12_q_net_x0,
    q_14 => delay13_q_net_x0,
    q_15 => delay14_q_net_x0,
    q_16 => delay15_q_net_x0
  );
  vector_delay1 : entity xil_defaultlib.psb3_0_vector_delay1_x0 
  port map (
    d_1 => slice0_y_net_x0,
    d_2 => slice1_y_net_x0,
    d_3 => slice2_y_net_x0,
    d_4 => slice3_y_net_x0,
    d_5 => slice4_y_net_x0,
    d_6 => slice5_y_net_x0,
    d_7 => slice6_y_net_x0,
    d_8 => slice7_y_net_x0,
    d_9 => slice8_y_net_x0,
    d_10 => slice9_y_net_x0,
    d_11 => slice10_y_net_x0,
    d_12 => slice11_y_net_x0,
    d_13 => slice12_y_net_x0,
    d_14 => slice13_y_net_x0,
    d_15 => slice14_y_net_x0,
    d_16 => slice15_y_net_x0,
    clk_1 => clk_net,
    ce_1 => ce_net,
    q_1 => delay0_q_net,
    q_2 => delay1_q_net,
    q_3 => delay2_q_net,
    q_4 => delay3_q_net,
    q_5 => delay4_q_net,
    q_6 => delay5_q_net,
    q_7 => delay6_q_net,
    q_8 => delay7_q_net,
    q_9 => delay8_q_net,
    q_10 => delay9_q_net,
    q_11 => delay10_q_net,
    q_12 => delay11_q_net,
    q_13 => delay12_q_net,
    q_14 => delay13_q_net,
    q_15 => delay14_q_net,
    q_16 => delay15_q_net
  );
  vector_slice : entity xil_defaultlib.psb3_0_vector_slice_x0 
  port map (
    in_1 => mult0_p_net,
    in_2 => mult1_p_net,
    in_3 => mult2_p_net,
    in_4 => mult3_p_net,
    in_5 => mult4_p_net,
    in_6 => mult5_p_net,
    in_7 => mult6_p_net,
    in_8 => mult7_p_net,
    in_9 => mult8_p_net,
    in_10 => mult9_p_net,
    in_11 => mult10_p_net,
    in_12 => mult11_p_net,
    in_13 => mult12_p_net,
    in_14 => mult13_p_net,
    in_15 => mult14_p_net,
    in_16 => mult15_p_net,
    out_1 => slice0_y_net_x1,
    out_2 => slice1_y_net_x1,
    out_3 => slice2_y_net_x1,
    out_4 => slice3_y_net_x1,
    out_5 => slice4_y_net_x1,
    out_6 => slice5_y_net_x1,
    out_7 => slice6_y_net_x1,
    out_8 => slice7_y_net_x1,
    out_9 => slice8_y_net_x1,
    out_10 => slice9_y_net_x1,
    out_11 => slice10_y_net_x1,
    out_12 => slice11_y_net_x1,
    out_13 => slice12_y_net_x1,
    out_14 => slice13_y_net_x1,
    out_15 => slice14_y_net_x1,
    out_16 => slice15_y_net_x1
  );
  vector_slice1 : entity xil_defaultlib.psb3_0_vector_slice1_x0 
  port map (
    in_1 => reinterpret0_output_port_net,
    in_2 => reinterpret1_output_port_net,
    in_3 => reinterpret2_output_port_net,
    in_4 => reinterpret3_output_port_net,
    in_5 => reinterpret4_output_port_net,
    in_6 => reinterpret5_output_port_net,
    in_7 => reinterpret6_output_port_net,
    in_8 => reinterpret7_output_port_net,
    in_9 => reinterpret8_output_port_net,
    in_10 => reinterpret9_output_port_net,
    in_11 => reinterpret10_output_port_net,
    in_12 => reinterpret11_output_port_net,
    in_13 => reinterpret12_output_port_net,
    in_14 => reinterpret13_output_port_net,
    in_15 => reinterpret14_output_port_net,
    in_16 => reinterpret15_output_port_net,
    out_1 => slice0_y_net_x0,
    out_2 => slice1_y_net_x0,
    out_3 => slice2_y_net_x0,
    out_4 => slice3_y_net_x0,
    out_5 => slice4_y_net_x0,
    out_6 => slice5_y_net_x0,
    out_7 => slice6_y_net_x0,
    out_8 => slice7_y_net_x0,
    out_9 => slice8_y_net_x0,
    out_10 => slice9_y_net_x0,
    out_11 => slice10_y_net_x0,
    out_12 => slice11_y_net_x0,
    out_13 => slice12_y_net_x0,
    out_14 => slice13_y_net_x0,
    out_15 => slice14_y_net_x0,
    out_16 => slice15_y_net_x0
  );
  vector_slice2 : entity xil_defaultlib.psb3_0_vector_slice2_x0 
  port map (
    in_1 => addsub0_s_net,
    in_2 => addsub1_s_net,
    in_3 => addsub2_s_net,
    in_4 => addsub3_s_net,
    in_5 => addsub4_s_net,
    in_6 => addsub5_s_net,
    in_7 => addsub6_s_net,
    in_8 => addsub7_s_net,
    in_9 => addsub8_s_net,
    in_10 => addsub9_s_net,
    in_11 => addsub10_s_net,
    in_12 => addsub11_s_net,
    in_13 => addsub12_s_net,
    in_14 => addsub13_s_net,
    in_15 => addsub14_s_net,
    in_16 => addsub15_s_net,
    out_1 => slice0_y_net,
    out_2 => slice1_y_net,
    out_3 => slice2_y_net,
    out_4 => slice3_y_net,
    out_5 => slice4_y_net,
    out_6 => slice5_y_net,
    out_7 => slice6_y_net,
    out_8 => slice7_y_net,
    out_9 => slice8_y_net,
    out_10 => slice9_y_net,
    out_11 => slice10_y_net,
    out_12 => slice11_y_net,
    out_13 => slice12_y_net,
    out_14 => slice13_y_net,
    out_15 => slice14_y_net,
    out_16 => slice15_y_net
  );
  vector_to_scalar : entity xil_defaultlib.psb3_0_vector_to_scalar_x0 
  port map (
    i_1 => delay0_q_net_x0,
    i_2 => delay1_q_net_x0,
    i_3 => delay2_q_net_x0,
    i_4 => delay3_q_net_x0,
    i_5 => delay4_q_net_x0,
    i_6 => delay5_q_net_x0,
    i_7 => delay6_q_net_x0,
    i_8 => delay7_q_net_x0,
    i_9 => delay8_q_net_x0,
    i_10 => delay9_q_net_x0,
    i_11 => delay10_q_net_x0,
    i_12 => delay11_q_net_x0,
    i_13 => delay12_q_net_x0,
    i_14 => delay13_q_net_x0,
    i_15 => delay14_q_net_x0,
    i_16 => delay15_q_net_x0,
    o => concat1_y_net_x1
  );
  vector_to_scalar1 : entity xil_defaultlib.psb3_0_vector_to_scalar1_x0 
  port map (
    i_1 => delay0_q_net,
    i_2 => delay1_q_net,
    i_3 => delay2_q_net,
    i_4 => delay3_q_net,
    i_5 => delay4_q_net,
    i_6 => delay5_q_net,
    i_7 => delay6_q_net,
    i_8 => delay7_q_net,
    i_9 => delay8_q_net,
    i_10 => delay9_q_net,
    i_11 => delay10_q_net,
    i_12 => delay11_q_net,
    i_13 => delay12_q_net,
    i_14 => delay13_q_net,
    i_15 => delay14_q_net,
    i_16 => delay15_q_net,
    o => concat1_y_net_x0
  );
  vector_to_scalar2 : entity xil_defaultlib.psb3_0_vector_to_scalar2_x1 
  port map (
    i_1 => slice0_y_net,
    i_2 => slice1_y_net,
    i_3 => slice2_y_net,
    i_4 => slice3_y_net,
    i_5 => slice4_y_net,
    i_6 => slice5_y_net,
    i_7 => slice6_y_net,
    i_8 => slice7_y_net,
    i_9 => slice8_y_net,
    i_10 => slice9_y_net,
    i_11 => slice10_y_net,
    i_12 => slice11_y_net,
    i_13 => slice12_y_net,
    i_14 => slice13_y_net,
    i_15 => slice14_y_net,
    i_16 => slice15_y_net,
    o => concat1_y_net
  );
  constant17 : entity xil_defaultlib.sysgen_constant_71e89d757c 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant17_op_net
  );
  convert : entity xil_defaultlib.psb3_0_xlconvert 
  generic map (
    bool_conversion => 1,
    din_arith => 1,
    din_bin_pt => 0,
    din_width => 1,
    dout_arith => 1,
    dout_bin_pt => 0,
    dout_width => 1,
    latency => 1,
    overflow => xlWrap,
    quantization => xlTruncate
  )
  port map (
    clr => '0',
    en => "1",
    din => expression_dout_net,
    clk => clk_net,
    ce => ce_net,
    dout => convert_dout_net
  );
  expression : entity xil_defaultlib.sysgen_expr_7c83532765 
  port map (
    clr => '0',
    a => concat1_y_net_x1,
    b => concat1_y_net_x0,
    s => concat1_y_net,
    clk => clk_net,
    ce => ce_net,
    dout => expression_dout_net
  );
  register_x0 : entity xil_defaultlib.psb3_0_xlregister 
  generic map (
    d_width => 1,
    init_value => b"0"
  )
  port map (
    d => constant17_op_net,
    rst => gin_tl_reset_net,
    en => convert_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => register_q_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Overflow Detector add_im_3/Vector Delay
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_delay_x1 is
  port (
    d_1 : in std_logic_vector( 1-1 downto 0 );
    d_2 : in std_logic_vector( 1-1 downto 0 );
    d_3 : in std_logic_vector( 1-1 downto 0 );
    d_4 : in std_logic_vector( 1-1 downto 0 );
    d_5 : in std_logic_vector( 1-1 downto 0 );
    d_6 : in std_logic_vector( 1-1 downto 0 );
    d_7 : in std_logic_vector( 1-1 downto 0 );
    d_8 : in std_logic_vector( 1-1 downto 0 );
    d_9 : in std_logic_vector( 1-1 downto 0 );
    d_10 : in std_logic_vector( 1-1 downto 0 );
    d_11 : in std_logic_vector( 1-1 downto 0 );
    d_12 : in std_logic_vector( 1-1 downto 0 );
    d_13 : in std_logic_vector( 1-1 downto 0 );
    d_14 : in std_logic_vector( 1-1 downto 0 );
    d_15 : in std_logic_vector( 1-1 downto 0 );
    d_16 : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    q_1 : out std_logic_vector( 1-1 downto 0 );
    q_2 : out std_logic_vector( 1-1 downto 0 );
    q_3 : out std_logic_vector( 1-1 downto 0 );
    q_4 : out std_logic_vector( 1-1 downto 0 );
    q_5 : out std_logic_vector( 1-1 downto 0 );
    q_6 : out std_logic_vector( 1-1 downto 0 );
    q_7 : out std_logic_vector( 1-1 downto 0 );
    q_8 : out std_logic_vector( 1-1 downto 0 );
    q_9 : out std_logic_vector( 1-1 downto 0 );
    q_10 : out std_logic_vector( 1-1 downto 0 );
    q_11 : out std_logic_vector( 1-1 downto 0 );
    q_12 : out std_logic_vector( 1-1 downto 0 );
    q_13 : out std_logic_vector( 1-1 downto 0 );
    q_14 : out std_logic_vector( 1-1 downto 0 );
    q_15 : out std_logic_vector( 1-1 downto 0 );
    q_16 : out std_logic_vector( 1-1 downto 0 )
  );
end psb3_0_vector_delay_x1;
architecture structural of psb3_0_vector_delay_x1 is 
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay0_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay11_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay12_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay10_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal delay13_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay7_q_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal slice9_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay9_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay14_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay15_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 1-1 downto 0 );
begin
  q_1 <= delay0_q_net;
  q_2 <= delay1_q_net;
  q_3 <= delay2_q_net;
  q_4 <= delay3_q_net;
  q_5 <= delay4_q_net;
  q_6 <= delay5_q_net;
  q_7 <= delay6_q_net;
  q_8 <= delay7_q_net;
  q_9 <= delay8_q_net;
  q_10 <= delay9_q_net;
  q_11 <= delay10_q_net;
  q_12 <= delay11_q_net;
  q_13 <= delay12_q_net;
  q_14 <= delay13_q_net;
  q_15 <= delay14_q_net;
  q_16 <= delay15_q_net;
  slice0_y_net <= d_1;
  slice1_y_net <= d_2;
  slice2_y_net <= d_3;
  slice3_y_net <= d_4;
  slice4_y_net <= d_5;
  slice5_y_net <= d_6;
  slice6_y_net <= d_7;
  slice7_y_net <= d_8;
  slice8_y_net <= d_9;
  slice9_y_net <= d_10;
  slice10_y_net <= d_11;
  slice11_y_net <= d_12;
  slice12_y_net <= d_13;
  slice13_y_net <= d_14;
  slice14_y_net <= d_15;
  slice15_y_net <= d_16;
  clk_net <= clk_1;
  ce_net <= ce_1;
  delay0 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice0_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay0_q_net
  );
  delay1 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice2_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay3 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice3_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  delay4 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice4_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net
  );
  delay5 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice5_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  delay6 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice6_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay6_q_net
  );
  delay7 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice7_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay7_q_net
  );
  delay8 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice8_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay8_q_net
  );
  delay9 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice9_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay9_q_net
  );
  delay10 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice10_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay10_q_net
  );
  delay11 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice11_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay11_q_net
  );
  delay12 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice12_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay12_q_net
  );
  delay13 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice13_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay13_q_net
  );
  delay14 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice14_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay14_q_net
  );
  delay15 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice15_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay15_q_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Overflow Detector add_im_3/Vector Delay1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_delay1_x1 is
  port (
    d_1 : in std_logic_vector( 1-1 downto 0 );
    d_2 : in std_logic_vector( 1-1 downto 0 );
    d_3 : in std_logic_vector( 1-1 downto 0 );
    d_4 : in std_logic_vector( 1-1 downto 0 );
    d_5 : in std_logic_vector( 1-1 downto 0 );
    d_6 : in std_logic_vector( 1-1 downto 0 );
    d_7 : in std_logic_vector( 1-1 downto 0 );
    d_8 : in std_logic_vector( 1-1 downto 0 );
    d_9 : in std_logic_vector( 1-1 downto 0 );
    d_10 : in std_logic_vector( 1-1 downto 0 );
    d_11 : in std_logic_vector( 1-1 downto 0 );
    d_12 : in std_logic_vector( 1-1 downto 0 );
    d_13 : in std_logic_vector( 1-1 downto 0 );
    d_14 : in std_logic_vector( 1-1 downto 0 );
    d_15 : in std_logic_vector( 1-1 downto 0 );
    d_16 : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    q_1 : out std_logic_vector( 1-1 downto 0 );
    q_2 : out std_logic_vector( 1-1 downto 0 );
    q_3 : out std_logic_vector( 1-1 downto 0 );
    q_4 : out std_logic_vector( 1-1 downto 0 );
    q_5 : out std_logic_vector( 1-1 downto 0 );
    q_6 : out std_logic_vector( 1-1 downto 0 );
    q_7 : out std_logic_vector( 1-1 downto 0 );
    q_8 : out std_logic_vector( 1-1 downto 0 );
    q_9 : out std_logic_vector( 1-1 downto 0 );
    q_10 : out std_logic_vector( 1-1 downto 0 );
    q_11 : out std_logic_vector( 1-1 downto 0 );
    q_12 : out std_logic_vector( 1-1 downto 0 );
    q_13 : out std_logic_vector( 1-1 downto 0 );
    q_14 : out std_logic_vector( 1-1 downto 0 );
    q_15 : out std_logic_vector( 1-1 downto 0 );
    q_16 : out std_logic_vector( 1-1 downto 0 )
  );
end psb3_0_vector_delay1_x1;
architecture structural of psb3_0_vector_delay1_x1 is 
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay11_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay12_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay0_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay10_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay13_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay14_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay15_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay7_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay9_q_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal slice1_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal slice9_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 1-1 downto 0 );
begin
  q_1 <= delay0_q_net;
  q_2 <= delay1_q_net;
  q_3 <= delay2_q_net;
  q_4 <= delay3_q_net;
  q_5 <= delay4_q_net;
  q_6 <= delay5_q_net;
  q_7 <= delay6_q_net;
  q_8 <= delay7_q_net;
  q_9 <= delay8_q_net;
  q_10 <= delay9_q_net;
  q_11 <= delay10_q_net;
  q_12 <= delay11_q_net;
  q_13 <= delay12_q_net;
  q_14 <= delay13_q_net;
  q_15 <= delay14_q_net;
  q_16 <= delay15_q_net;
  slice0_y_net <= d_1;
  slice1_y_net <= d_2;
  slice2_y_net <= d_3;
  slice3_y_net <= d_4;
  slice4_y_net <= d_5;
  slice5_y_net <= d_6;
  slice6_y_net <= d_7;
  slice7_y_net <= d_8;
  slice8_y_net <= d_9;
  slice9_y_net <= d_10;
  slice10_y_net <= d_11;
  slice11_y_net <= d_12;
  slice12_y_net <= d_13;
  slice13_y_net <= d_14;
  slice14_y_net <= d_15;
  slice15_y_net <= d_16;
  clk_net <= clk_1;
  ce_net <= ce_1;
  delay0 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice0_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay0_q_net
  );
  delay1 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice2_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay3 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice3_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  delay4 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice4_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net
  );
  delay5 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice5_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  delay6 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice6_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay6_q_net
  );
  delay7 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice7_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay7_q_net
  );
  delay8 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice8_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay8_q_net
  );
  delay9 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice9_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay9_q_net
  );
  delay10 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice10_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay10_q_net
  );
  delay11 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice11_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay11_q_net
  );
  delay12 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice12_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay12_q_net
  );
  delay13 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice13_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay13_q_net
  );
  delay14 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice14_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay14_q_net
  );
  delay15 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice15_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay15_q_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Overflow Detector add_im_3/Vector Slice
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_slice_x1 is
  port (
    in_1 : in std_logic_vector( 16-1 downto 0 );
    in_2 : in std_logic_vector( 16-1 downto 0 );
    in_3 : in std_logic_vector( 16-1 downto 0 );
    in_4 : in std_logic_vector( 16-1 downto 0 );
    in_5 : in std_logic_vector( 16-1 downto 0 );
    in_6 : in std_logic_vector( 16-1 downto 0 );
    in_7 : in std_logic_vector( 16-1 downto 0 );
    in_8 : in std_logic_vector( 16-1 downto 0 );
    in_9 : in std_logic_vector( 16-1 downto 0 );
    in_10 : in std_logic_vector( 16-1 downto 0 );
    in_11 : in std_logic_vector( 16-1 downto 0 );
    in_12 : in std_logic_vector( 16-1 downto 0 );
    in_13 : in std_logic_vector( 16-1 downto 0 );
    in_14 : in std_logic_vector( 16-1 downto 0 );
    in_15 : in std_logic_vector( 16-1 downto 0 );
    in_16 : in std_logic_vector( 16-1 downto 0 );
    out_1 : out std_logic_vector( 1-1 downto 0 );
    out_2 : out std_logic_vector( 1-1 downto 0 );
    out_3 : out std_logic_vector( 1-1 downto 0 );
    out_4 : out std_logic_vector( 1-1 downto 0 );
    out_5 : out std_logic_vector( 1-1 downto 0 );
    out_6 : out std_logic_vector( 1-1 downto 0 );
    out_7 : out std_logic_vector( 1-1 downto 0 );
    out_8 : out std_logic_vector( 1-1 downto 0 );
    out_9 : out std_logic_vector( 1-1 downto 0 );
    out_10 : out std_logic_vector( 1-1 downto 0 );
    out_11 : out std_logic_vector( 1-1 downto 0 );
    out_12 : out std_logic_vector( 1-1 downto 0 );
    out_13 : out std_logic_vector( 1-1 downto 0 );
    out_14 : out std_logic_vector( 1-1 downto 0 );
    out_15 : out std_logic_vector( 1-1 downto 0 );
    out_16 : out std_logic_vector( 1-1 downto 0 )
  );
end psb3_0_vector_slice_x1;
architecture structural of psb3_0_vector_slice_x1 is 
  signal slice4_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 1-1 downto 0 );
  signal mult0_p_net : std_logic_vector( 16-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 1-1 downto 0 );
  signal mult3_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult4_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult8_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult5_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult6_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult1_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult13_p_net : std_logic_vector( 16-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 1-1 downto 0 );
  signal mult11_p_net : std_logic_vector( 16-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 1-1 downto 0 );
  signal mult2_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult7_p_net : std_logic_vector( 16-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 1-1 downto 0 );
  signal mult9_p_net : std_logic_vector( 16-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 1-1 downto 0 );
  signal mult10_p_net : std_logic_vector( 16-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 1-1 downto 0 );
  signal mult12_p_net : std_logic_vector( 16-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 1-1 downto 0 );
  signal mult14_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult15_p_net : std_logic_vector( 16-1 downto 0 );
begin
  out_1 <= slice0_y_net;
  out_2 <= slice1_y_net;
  out_3 <= slice2_y_net;
  out_4 <= slice3_y_net;
  out_5 <= slice4_y_net;
  out_6 <= slice5_y_net;
  out_7 <= slice6_y_net;
  out_8 <= slice7_y_net;
  out_9 <= slice8_y_net;
  out_10 <= slice9_y_net;
  out_11 <= slice10_y_net;
  out_12 <= slice11_y_net;
  out_13 <= slice12_y_net;
  out_14 <= slice13_y_net;
  out_15 <= slice14_y_net;
  out_16 <= slice15_y_net;
  mult0_p_net <= in_1;
  mult1_p_net <= in_2;
  mult2_p_net <= in_3;
  mult3_p_net <= in_4;
  mult4_p_net <= in_5;
  mult5_p_net <= in_6;
  mult6_p_net <= in_7;
  mult7_p_net <= in_8;
  mult8_p_net <= in_9;
  mult9_p_net <= in_10;
  mult10_p_net <= in_11;
  mult11_p_net <= in_12;
  mult12_p_net <= in_13;
  mult13_p_net <= in_14;
  mult14_p_net <= in_15;
  mult15_p_net <= in_16;
  slice0 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult0_p_net,
    y => slice0_y_net
  );
  slice1 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult1_p_net,
    y => slice1_y_net
  );
  slice2 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult2_p_net,
    y => slice2_y_net
  );
  slice3 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult3_p_net,
    y => slice3_y_net
  );
  slice4 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult4_p_net,
    y => slice4_y_net
  );
  slice5 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult5_p_net,
    y => slice5_y_net
  );
  slice6 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult6_p_net,
    y => slice6_y_net
  );
  slice7 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult7_p_net,
    y => slice7_y_net
  );
  slice8 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult8_p_net,
    y => slice8_y_net
  );
  slice9 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult9_p_net,
    y => slice9_y_net
  );
  slice10 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult10_p_net,
    y => slice10_y_net
  );
  slice11 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult11_p_net,
    y => slice11_y_net
  );
  slice12 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult12_p_net,
    y => slice12_y_net
  );
  slice13 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult13_p_net,
    y => slice13_y_net
  );
  slice14 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult14_p_net,
    y => slice14_y_net
  );
  slice15 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult15_p_net,
    y => slice15_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Overflow Detector add_im_3/Vector Slice1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_slice1_x1 is
  port (
    in_1 : in std_logic_vector( 16-1 downto 0 );
    in_2 : in std_logic_vector( 16-1 downto 0 );
    in_3 : in std_logic_vector( 16-1 downto 0 );
    in_4 : in std_logic_vector( 16-1 downto 0 );
    in_5 : in std_logic_vector( 16-1 downto 0 );
    in_6 : in std_logic_vector( 16-1 downto 0 );
    in_7 : in std_logic_vector( 16-1 downto 0 );
    in_8 : in std_logic_vector( 16-1 downto 0 );
    in_9 : in std_logic_vector( 16-1 downto 0 );
    in_10 : in std_logic_vector( 16-1 downto 0 );
    in_11 : in std_logic_vector( 16-1 downto 0 );
    in_12 : in std_logic_vector( 16-1 downto 0 );
    in_13 : in std_logic_vector( 16-1 downto 0 );
    in_14 : in std_logic_vector( 16-1 downto 0 );
    in_15 : in std_logic_vector( 16-1 downto 0 );
    in_16 : in std_logic_vector( 16-1 downto 0 );
    out_1 : out std_logic_vector( 1-1 downto 0 );
    out_2 : out std_logic_vector( 1-1 downto 0 );
    out_3 : out std_logic_vector( 1-1 downto 0 );
    out_4 : out std_logic_vector( 1-1 downto 0 );
    out_5 : out std_logic_vector( 1-1 downto 0 );
    out_6 : out std_logic_vector( 1-1 downto 0 );
    out_7 : out std_logic_vector( 1-1 downto 0 );
    out_8 : out std_logic_vector( 1-1 downto 0 );
    out_9 : out std_logic_vector( 1-1 downto 0 );
    out_10 : out std_logic_vector( 1-1 downto 0 );
    out_11 : out std_logic_vector( 1-1 downto 0 );
    out_12 : out std_logic_vector( 1-1 downto 0 );
    out_13 : out std_logic_vector( 1-1 downto 0 );
    out_14 : out std_logic_vector( 1-1 downto 0 );
    out_15 : out std_logic_vector( 1-1 downto 0 );
    out_16 : out std_logic_vector( 1-1 downto 0 )
  );
end psb3_0_vector_slice1_x1;
architecture structural of psb3_0_vector_slice1_x1 is 
  signal slice1_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
begin
  out_1 <= slice0_y_net;
  out_2 <= slice1_y_net;
  out_3 <= slice2_y_net;
  out_4 <= slice3_y_net;
  out_5 <= slice4_y_net;
  out_6 <= slice5_y_net;
  out_7 <= slice6_y_net;
  out_8 <= slice7_y_net;
  out_9 <= slice8_y_net;
  out_10 <= slice9_y_net;
  out_11 <= slice10_y_net;
  out_12 <= slice11_y_net;
  out_13 <= slice12_y_net;
  out_14 <= slice13_y_net;
  out_15 <= slice14_y_net;
  out_16 <= slice15_y_net;
  reinterpret0_output_port_net <= in_1;
  reinterpret1_output_port_net <= in_2;
  reinterpret2_output_port_net <= in_3;
  reinterpret3_output_port_net <= in_4;
  reinterpret4_output_port_net <= in_5;
  reinterpret5_output_port_net <= in_6;
  reinterpret6_output_port_net <= in_7;
  reinterpret7_output_port_net <= in_8;
  reinterpret8_output_port_net <= in_9;
  reinterpret9_output_port_net <= in_10;
  reinterpret10_output_port_net <= in_11;
  reinterpret11_output_port_net <= in_12;
  reinterpret12_output_port_net <= in_13;
  reinterpret13_output_port_net <= in_14;
  reinterpret14_output_port_net <= in_15;
  reinterpret15_output_port_net <= in_16;
  slice0 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret0_output_port_net,
    y => slice0_y_net
  );
  slice1 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret1_output_port_net,
    y => slice1_y_net
  );
  slice2 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret2_output_port_net,
    y => slice2_y_net
  );
  slice3 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret3_output_port_net,
    y => slice3_y_net
  );
  slice4 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret4_output_port_net,
    y => slice4_y_net
  );
  slice5 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret5_output_port_net,
    y => slice5_y_net
  );
  slice6 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret6_output_port_net,
    y => slice6_y_net
  );
  slice7 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret7_output_port_net,
    y => slice7_y_net
  );
  slice8 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret8_output_port_net,
    y => slice8_y_net
  );
  slice9 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret9_output_port_net,
    y => slice9_y_net
  );
  slice10 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret10_output_port_net,
    y => slice10_y_net
  );
  slice11 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret11_output_port_net,
    y => slice11_y_net
  );
  slice12 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret12_output_port_net,
    y => slice12_y_net
  );
  slice13 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret13_output_port_net,
    y => slice13_y_net
  );
  slice14 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret14_output_port_net,
    y => slice14_y_net
  );
  slice15 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret15_output_port_net,
    y => slice15_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Overflow Detector add_im_3/Vector Slice2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_slice2_x1 is
  port (
    in_1 : in std_logic_vector( 16-1 downto 0 );
    in_2 : in std_logic_vector( 16-1 downto 0 );
    in_3 : in std_logic_vector( 16-1 downto 0 );
    in_4 : in std_logic_vector( 16-1 downto 0 );
    in_5 : in std_logic_vector( 16-1 downto 0 );
    in_6 : in std_logic_vector( 16-1 downto 0 );
    in_7 : in std_logic_vector( 16-1 downto 0 );
    in_8 : in std_logic_vector( 16-1 downto 0 );
    in_9 : in std_logic_vector( 16-1 downto 0 );
    in_10 : in std_logic_vector( 16-1 downto 0 );
    in_11 : in std_logic_vector( 16-1 downto 0 );
    in_12 : in std_logic_vector( 16-1 downto 0 );
    in_13 : in std_logic_vector( 16-1 downto 0 );
    in_14 : in std_logic_vector( 16-1 downto 0 );
    in_15 : in std_logic_vector( 16-1 downto 0 );
    in_16 : in std_logic_vector( 16-1 downto 0 );
    out_1 : out std_logic_vector( 1-1 downto 0 );
    out_2 : out std_logic_vector( 1-1 downto 0 );
    out_3 : out std_logic_vector( 1-1 downto 0 );
    out_4 : out std_logic_vector( 1-1 downto 0 );
    out_5 : out std_logic_vector( 1-1 downto 0 );
    out_6 : out std_logic_vector( 1-1 downto 0 );
    out_7 : out std_logic_vector( 1-1 downto 0 );
    out_8 : out std_logic_vector( 1-1 downto 0 );
    out_9 : out std_logic_vector( 1-1 downto 0 );
    out_10 : out std_logic_vector( 1-1 downto 0 );
    out_11 : out std_logic_vector( 1-1 downto 0 );
    out_12 : out std_logic_vector( 1-1 downto 0 );
    out_13 : out std_logic_vector( 1-1 downto 0 );
    out_14 : out std_logic_vector( 1-1 downto 0 );
    out_15 : out std_logic_vector( 1-1 downto 0 );
    out_16 : out std_logic_vector( 1-1 downto 0 )
  );
end psb3_0_vector_slice2_x1;
architecture structural of psb3_0_vector_slice2_x1 is 
  signal slice2_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 1-1 downto 0 );
  signal addsub0_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub3_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub8_s_net : std_logic_vector( 16-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 1-1 downto 0 );
  signal addsub7_s_net : std_logic_vector( 16-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 1-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub10_s_net : std_logic_vector( 16-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 1-1 downto 0 );
  signal addsub11_s_net : std_logic_vector( 16-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 1-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub5_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub6_s_net : std_logic_vector( 16-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 1-1 downto 0 );
  signal addsub9_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub12_s_net : std_logic_vector( 16-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 1-1 downto 0 );
  signal addsub15_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub13_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub14_s_net : std_logic_vector( 16-1 downto 0 );
begin
  out_1 <= slice0_y_net;
  out_2 <= slice1_y_net;
  out_3 <= slice2_y_net;
  out_4 <= slice3_y_net;
  out_5 <= slice4_y_net;
  out_6 <= slice5_y_net;
  out_7 <= slice6_y_net;
  out_8 <= slice7_y_net;
  out_9 <= slice8_y_net;
  out_10 <= slice9_y_net;
  out_11 <= slice10_y_net;
  out_12 <= slice11_y_net;
  out_13 <= slice12_y_net;
  out_14 <= slice13_y_net;
  out_15 <= slice14_y_net;
  out_16 <= slice15_y_net;
  addsub0_s_net <= in_1;
  addsub1_s_net <= in_2;
  addsub2_s_net <= in_3;
  addsub3_s_net <= in_4;
  addsub4_s_net <= in_5;
  addsub5_s_net <= in_6;
  addsub6_s_net <= in_7;
  addsub7_s_net <= in_8;
  addsub8_s_net <= in_9;
  addsub9_s_net <= in_10;
  addsub10_s_net <= in_11;
  addsub11_s_net <= in_12;
  addsub12_s_net <= in_13;
  addsub13_s_net <= in_14;
  addsub14_s_net <= in_15;
  addsub15_s_net <= in_16;
  slice0 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub0_s_net,
    y => slice0_y_net
  );
  slice1 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub1_s_net,
    y => slice1_y_net
  );
  slice2 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub2_s_net,
    y => slice2_y_net
  );
  slice3 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub3_s_net,
    y => slice3_y_net
  );
  slice4 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub4_s_net,
    y => slice4_y_net
  );
  slice5 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub5_s_net,
    y => slice5_y_net
  );
  slice6 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub6_s_net,
    y => slice6_y_net
  );
  slice7 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub7_s_net,
    y => slice7_y_net
  );
  slice8 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub8_s_net,
    y => slice8_y_net
  );
  slice9 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub9_s_net,
    y => slice9_y_net
  );
  slice10 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub10_s_net,
    y => slice10_y_net
  );
  slice11 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub11_s_net,
    y => slice11_y_net
  );
  slice12 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub12_s_net,
    y => slice12_y_net
  );
  slice13 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub13_s_net,
    y => slice13_y_net
  );
  slice14 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub14_s_net,
    y => slice14_y_net
  );
  slice15 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub15_s_net,
    y => slice15_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Overflow Detector add_im_3/Vector to Scalar
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_to_scalar_x1 is
  port (
    i_1 : in std_logic_vector( 1-1 downto 0 );
    i_2 : in std_logic_vector( 1-1 downto 0 );
    i_3 : in std_logic_vector( 1-1 downto 0 );
    i_4 : in std_logic_vector( 1-1 downto 0 );
    i_5 : in std_logic_vector( 1-1 downto 0 );
    i_6 : in std_logic_vector( 1-1 downto 0 );
    i_7 : in std_logic_vector( 1-1 downto 0 );
    i_8 : in std_logic_vector( 1-1 downto 0 );
    i_9 : in std_logic_vector( 1-1 downto 0 );
    i_10 : in std_logic_vector( 1-1 downto 0 );
    i_11 : in std_logic_vector( 1-1 downto 0 );
    i_12 : in std_logic_vector( 1-1 downto 0 );
    i_13 : in std_logic_vector( 1-1 downto 0 );
    i_14 : in std_logic_vector( 1-1 downto 0 );
    i_15 : in std_logic_vector( 1-1 downto 0 );
    i_16 : in std_logic_vector( 1-1 downto 0 );
    o : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_vector_to_scalar_x1;
architecture structural of psb3_0_vector_to_scalar_x1 is 
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay0_q_net : std_logic_vector( 1-1 downto 0 );
  signal concat1_y_net : std_logic_vector( 16-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay11_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay7_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay9_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay10_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay15_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay13_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay12_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay14_q_net : std_logic_vector( 1-1 downto 0 );
begin
  o <= concat1_y_net;
  delay0_q_net <= i_1;
  delay1_q_net <= i_2;
  delay2_q_net <= i_3;
  delay3_q_net <= i_4;
  delay4_q_net <= i_5;
  delay5_q_net <= i_6;
  delay6_q_net <= i_7;
  delay7_q_net <= i_8;
  delay8_q_net <= i_9;
  delay9_q_net <= i_10;
  delay10_q_net <= i_11;
  delay11_q_net <= i_12;
  delay12_q_net <= i_13;
  delay13_q_net <= i_14;
  delay14_q_net <= i_15;
  delay15_q_net <= i_16;
  concat1 : entity xil_defaultlib.sysgen_concat_d977c66e35 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => delay15_q_net,
    in1 => delay14_q_net,
    in2 => delay13_q_net,
    in3 => delay12_q_net,
    in4 => delay11_q_net,
    in5 => delay10_q_net,
    in6 => delay9_q_net,
    in7 => delay8_q_net,
    in8 => delay7_q_net,
    in9 => delay6_q_net,
    in10 => delay5_q_net,
    in11 => delay4_q_net,
    in12 => delay3_q_net,
    in13 => delay2_q_net,
    in14 => delay1_q_net,
    in15 => delay0_q_net,
    y => concat1_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Overflow Detector add_im_3/Vector to Scalar1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_to_scalar1_x1 is
  port (
    i_1 : in std_logic_vector( 1-1 downto 0 );
    i_2 : in std_logic_vector( 1-1 downto 0 );
    i_3 : in std_logic_vector( 1-1 downto 0 );
    i_4 : in std_logic_vector( 1-1 downto 0 );
    i_5 : in std_logic_vector( 1-1 downto 0 );
    i_6 : in std_logic_vector( 1-1 downto 0 );
    i_7 : in std_logic_vector( 1-1 downto 0 );
    i_8 : in std_logic_vector( 1-1 downto 0 );
    i_9 : in std_logic_vector( 1-1 downto 0 );
    i_10 : in std_logic_vector( 1-1 downto 0 );
    i_11 : in std_logic_vector( 1-1 downto 0 );
    i_12 : in std_logic_vector( 1-1 downto 0 );
    i_13 : in std_logic_vector( 1-1 downto 0 );
    i_14 : in std_logic_vector( 1-1 downto 0 );
    i_15 : in std_logic_vector( 1-1 downto 0 );
    i_16 : in std_logic_vector( 1-1 downto 0 );
    o : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_vector_to_scalar1_x1;
architecture structural of psb3_0_vector_to_scalar1_x1 is 
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay0_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay11_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay12_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay10_q_net : std_logic_vector( 1-1 downto 0 );
  signal concat1_y_net : std_logic_vector( 16-1 downto 0 );
  signal delay9_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay15_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay13_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay7_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay14_q_net : std_logic_vector( 1-1 downto 0 );
begin
  o <= concat1_y_net;
  delay0_q_net <= i_1;
  delay1_q_net <= i_2;
  delay2_q_net <= i_3;
  delay3_q_net <= i_4;
  delay4_q_net <= i_5;
  delay5_q_net <= i_6;
  delay6_q_net <= i_7;
  delay7_q_net <= i_8;
  delay8_q_net <= i_9;
  delay9_q_net <= i_10;
  delay10_q_net <= i_11;
  delay11_q_net <= i_12;
  delay12_q_net <= i_13;
  delay13_q_net <= i_14;
  delay14_q_net <= i_15;
  delay15_q_net <= i_16;
  concat1 : entity xil_defaultlib.sysgen_concat_d977c66e35 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => delay15_q_net,
    in1 => delay14_q_net,
    in2 => delay13_q_net,
    in3 => delay12_q_net,
    in4 => delay11_q_net,
    in5 => delay10_q_net,
    in6 => delay9_q_net,
    in7 => delay8_q_net,
    in8 => delay7_q_net,
    in9 => delay6_q_net,
    in10 => delay5_q_net,
    in11 => delay4_q_net,
    in12 => delay3_q_net,
    in13 => delay2_q_net,
    in14 => delay1_q_net,
    in15 => delay0_q_net,
    y => concat1_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Overflow Detector add_im_3/Vector to Scalar2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_to_scalar2 is
  port (
    i_1 : in std_logic_vector( 1-1 downto 0 );
    i_2 : in std_logic_vector( 1-1 downto 0 );
    i_3 : in std_logic_vector( 1-1 downto 0 );
    i_4 : in std_logic_vector( 1-1 downto 0 );
    i_5 : in std_logic_vector( 1-1 downto 0 );
    i_6 : in std_logic_vector( 1-1 downto 0 );
    i_7 : in std_logic_vector( 1-1 downto 0 );
    i_8 : in std_logic_vector( 1-1 downto 0 );
    i_9 : in std_logic_vector( 1-1 downto 0 );
    i_10 : in std_logic_vector( 1-1 downto 0 );
    i_11 : in std_logic_vector( 1-1 downto 0 );
    i_12 : in std_logic_vector( 1-1 downto 0 );
    i_13 : in std_logic_vector( 1-1 downto 0 );
    i_14 : in std_logic_vector( 1-1 downto 0 );
    i_15 : in std_logic_vector( 1-1 downto 0 );
    i_16 : in std_logic_vector( 1-1 downto 0 );
    o : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_vector_to_scalar2;
architecture structural of psb3_0_vector_to_scalar2 is 
  signal slice7_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 1-1 downto 0 );
  signal concat1_y_net : std_logic_vector( 16-1 downto 0 );
begin
  o <= concat1_y_net;
  slice0_y_net <= i_1;
  slice1_y_net <= i_2;
  slice2_y_net <= i_3;
  slice3_y_net <= i_4;
  slice4_y_net <= i_5;
  slice5_y_net <= i_6;
  slice6_y_net <= i_7;
  slice7_y_net <= i_8;
  slice8_y_net <= i_9;
  slice9_y_net <= i_10;
  slice10_y_net <= i_11;
  slice11_y_net <= i_12;
  slice12_y_net <= i_13;
  slice13_y_net <= i_14;
  slice14_y_net <= i_15;
  slice15_y_net <= i_16;
  concat1 : entity xil_defaultlib.sysgen_concat_d977c66e35 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => slice15_y_net,
    in1 => slice14_y_net,
    in2 => slice13_y_net,
    in3 => slice12_y_net,
    in4 => slice11_y_net,
    in5 => slice10_y_net,
    in6 => slice9_y_net,
    in7 => slice8_y_net,
    in8 => slice7_y_net,
    in9 => slice6_y_net,
    in10 => slice5_y_net,
    in11 => slice4_y_net,
    in12 => slice3_y_net,
    in13 => slice2_y_net,
    in14 => slice1_y_net,
    in15 => slice0_y_net,
    y => concat1_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Overflow Detector add_im_3
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_overflow_detector_add_im_3 is
  port (
    rst : in std_logic_vector( 1-1 downto 0 );
    a_1 : in std_logic_vector( 16-1 downto 0 );
    b_1 : in std_logic_vector( 16-1 downto 0 );
    s_1 : in std_logic_vector( 16-1 downto 0 );
    a_2 : in std_logic_vector( 16-1 downto 0 );
    a_3 : in std_logic_vector( 16-1 downto 0 );
    a_4 : in std_logic_vector( 16-1 downto 0 );
    a_5 : in std_logic_vector( 16-1 downto 0 );
    a_6 : in std_logic_vector( 16-1 downto 0 );
    a_7 : in std_logic_vector( 16-1 downto 0 );
    a_8 : in std_logic_vector( 16-1 downto 0 );
    a_9 : in std_logic_vector( 16-1 downto 0 );
    a_10 : in std_logic_vector( 16-1 downto 0 );
    a_11 : in std_logic_vector( 16-1 downto 0 );
    a_12 : in std_logic_vector( 16-1 downto 0 );
    a_13 : in std_logic_vector( 16-1 downto 0 );
    a_14 : in std_logic_vector( 16-1 downto 0 );
    a_15 : in std_logic_vector( 16-1 downto 0 );
    a_16 : in std_logic_vector( 16-1 downto 0 );
    b_2 : in std_logic_vector( 16-1 downto 0 );
    b_3 : in std_logic_vector( 16-1 downto 0 );
    b_4 : in std_logic_vector( 16-1 downto 0 );
    b_5 : in std_logic_vector( 16-1 downto 0 );
    b_6 : in std_logic_vector( 16-1 downto 0 );
    b_7 : in std_logic_vector( 16-1 downto 0 );
    b_8 : in std_logic_vector( 16-1 downto 0 );
    b_9 : in std_logic_vector( 16-1 downto 0 );
    b_10 : in std_logic_vector( 16-1 downto 0 );
    b_11 : in std_logic_vector( 16-1 downto 0 );
    b_12 : in std_logic_vector( 16-1 downto 0 );
    b_13 : in std_logic_vector( 16-1 downto 0 );
    b_14 : in std_logic_vector( 16-1 downto 0 );
    b_15 : in std_logic_vector( 16-1 downto 0 );
    b_16 : in std_logic_vector( 16-1 downto 0 );
    s_2 : in std_logic_vector( 16-1 downto 0 );
    s_3 : in std_logic_vector( 16-1 downto 0 );
    s_4 : in std_logic_vector( 16-1 downto 0 );
    s_5 : in std_logic_vector( 16-1 downto 0 );
    s_6 : in std_logic_vector( 16-1 downto 0 );
    s_7 : in std_logic_vector( 16-1 downto 0 );
    s_8 : in std_logic_vector( 16-1 downto 0 );
    s_9 : in std_logic_vector( 16-1 downto 0 );
    s_10 : in std_logic_vector( 16-1 downto 0 );
    s_11 : in std_logic_vector( 16-1 downto 0 );
    s_12 : in std_logic_vector( 16-1 downto 0 );
    s_13 : in std_logic_vector( 16-1 downto 0 );
    s_14 : in std_logic_vector( 16-1 downto 0 );
    s_15 : in std_logic_vector( 16-1 downto 0 );
    s_16 : in std_logic_vector( 16-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    ov : out std_logic_vector( 1-1 downto 0 )
  );
end psb3_0_overflow_detector_add_im_3;
architecture structural of psb3_0_overflow_detector_add_im_3 is 
  signal mult14_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub0_s_net : std_logic_vector( 16-1 downto 0 );
  signal gin_tl_reset_net : std_logic_vector( 1-1 downto 0 );
  signal mult5_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult12_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mult15_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mult7_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult9_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult8_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult11_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult13_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult2_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult4_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult0_p_net : std_logic_vector( 16-1 downto 0 );
  signal register_q_net : std_logic_vector( 1-1 downto 0 );
  signal mult1_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult3_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult6_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult10_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub8_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub11_s_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub6_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub5_s_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub12_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub3_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub14_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub15_s_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub7_s_net : std_logic_vector( 16-1 downto 0 );
  signal ce_net : std_logic;
  signal delay2_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal delay3_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal addsub9_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub10_s_net : std_logic_vector( 16-1 downto 0 );
  signal delay0_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal addsub13_s_net : std_logic_vector( 16-1 downto 0 );
  signal delay4_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay5_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay6_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay8_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal delay7_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay9_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay10_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice14_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal slice6_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal delay0_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice11_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay12_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay13_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice14_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice1_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice15_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice15_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice9_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice2_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice5_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal delay7_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice13_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal slice13_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice4_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay14_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay11_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice8_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal slice6_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice7_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice10_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay12_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay15_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice12_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice3_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal delay15_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice5_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay9_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice8_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice11_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal slice7_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal slice0_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal delay13_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice3_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice12_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal delay14_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice9_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal slice4_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay10_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay11_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice0_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice1_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice2_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice10_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal concat1_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 1-1 downto 0 );
  signal constant17_op_net : std_logic_vector( 1-1 downto 0 );
  signal expression_dout_net : std_logic_vector( 1-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 1-1 downto 0 );
  signal concat1_y_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal concat1_y_net_x1 : std_logic_vector( 16-1 downto 0 );
  signal convert_dout_net : std_logic_vector( 1-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 1-1 downto 0 );
begin
  ov <= register_q_net;
  gin_tl_reset_net <= rst;
  mult0_p_net <= a_1;
  reinterpret0_output_port_net <= b_1;
  addsub0_s_net <= s_1;
  mult1_p_net <= a_2;
  mult2_p_net <= a_3;
  mult3_p_net <= a_4;
  mult4_p_net <= a_5;
  mult5_p_net <= a_6;
  mult6_p_net <= a_7;
  mult7_p_net <= a_8;
  mult8_p_net <= a_9;
  mult9_p_net <= a_10;
  mult10_p_net <= a_11;
  mult11_p_net <= a_12;
  mult12_p_net <= a_13;
  mult13_p_net <= a_14;
  mult14_p_net <= a_15;
  mult15_p_net <= a_16;
  reinterpret1_output_port_net <= b_2;
  reinterpret2_output_port_net <= b_3;
  reinterpret3_output_port_net <= b_4;
  reinterpret4_output_port_net <= b_5;
  reinterpret5_output_port_net <= b_6;
  reinterpret6_output_port_net <= b_7;
  reinterpret7_output_port_net <= b_8;
  reinterpret8_output_port_net <= b_9;
  reinterpret9_output_port_net <= b_10;
  reinterpret10_output_port_net <= b_11;
  reinterpret11_output_port_net <= b_12;
  reinterpret12_output_port_net <= b_13;
  reinterpret13_output_port_net <= b_14;
  reinterpret14_output_port_net <= b_15;
  reinterpret15_output_port_net <= b_16;
  addsub1_s_net <= s_2;
  addsub2_s_net <= s_3;
  addsub3_s_net <= s_4;
  addsub4_s_net <= s_5;
  addsub5_s_net <= s_6;
  addsub6_s_net <= s_7;
  addsub7_s_net <= s_8;
  addsub8_s_net <= s_9;
  addsub9_s_net <= s_10;
  addsub10_s_net <= s_11;
  addsub11_s_net <= s_12;
  addsub12_s_net <= s_13;
  addsub13_s_net <= s_14;
  addsub14_s_net <= s_15;
  addsub15_s_net <= s_16;
  clk_net <= clk_1;
  ce_net <= ce_1;
  vector_delay : entity xil_defaultlib.psb3_0_vector_delay_x1 
  port map (
    d_1 => slice0_y_net_x1,
    d_2 => slice1_y_net_x1,
    d_3 => slice2_y_net_x1,
    d_4 => slice3_y_net_x1,
    d_5 => slice4_y_net_x1,
    d_6 => slice5_y_net_x1,
    d_7 => slice6_y_net_x1,
    d_8 => slice7_y_net_x1,
    d_9 => slice8_y_net_x1,
    d_10 => slice9_y_net_x1,
    d_11 => slice10_y_net_x1,
    d_12 => slice11_y_net_x1,
    d_13 => slice12_y_net_x1,
    d_14 => slice13_y_net_x1,
    d_15 => slice14_y_net_x1,
    d_16 => slice15_y_net_x1,
    clk_1 => clk_net,
    ce_1 => ce_net,
    q_1 => delay0_q_net_x0,
    q_2 => delay1_q_net_x0,
    q_3 => delay2_q_net_x0,
    q_4 => delay3_q_net_x0,
    q_5 => delay4_q_net_x0,
    q_6 => delay5_q_net_x0,
    q_7 => delay6_q_net_x0,
    q_8 => delay7_q_net_x0,
    q_9 => delay8_q_net_x0,
    q_10 => delay9_q_net_x0,
    q_11 => delay10_q_net_x0,
    q_12 => delay11_q_net_x0,
    q_13 => delay12_q_net_x0,
    q_14 => delay13_q_net_x0,
    q_15 => delay14_q_net_x0,
    q_16 => delay15_q_net_x0
  );
  vector_delay1 : entity xil_defaultlib.psb3_0_vector_delay1_x1 
  port map (
    d_1 => slice0_y_net_x0,
    d_2 => slice1_y_net_x0,
    d_3 => slice2_y_net_x0,
    d_4 => slice3_y_net_x0,
    d_5 => slice4_y_net_x0,
    d_6 => slice5_y_net_x0,
    d_7 => slice6_y_net_x0,
    d_8 => slice7_y_net_x0,
    d_9 => slice8_y_net_x0,
    d_10 => slice9_y_net_x0,
    d_11 => slice10_y_net_x0,
    d_12 => slice11_y_net_x0,
    d_13 => slice12_y_net_x0,
    d_14 => slice13_y_net_x0,
    d_15 => slice14_y_net_x0,
    d_16 => slice15_y_net_x0,
    clk_1 => clk_net,
    ce_1 => ce_net,
    q_1 => delay0_q_net,
    q_2 => delay1_q_net,
    q_3 => delay2_q_net,
    q_4 => delay3_q_net,
    q_5 => delay4_q_net,
    q_6 => delay5_q_net,
    q_7 => delay6_q_net,
    q_8 => delay7_q_net,
    q_9 => delay8_q_net,
    q_10 => delay9_q_net,
    q_11 => delay10_q_net,
    q_12 => delay11_q_net,
    q_13 => delay12_q_net,
    q_14 => delay13_q_net,
    q_15 => delay14_q_net,
    q_16 => delay15_q_net
  );
  vector_slice : entity xil_defaultlib.psb3_0_vector_slice_x1 
  port map (
    in_1 => mult0_p_net,
    in_2 => mult1_p_net,
    in_3 => mult2_p_net,
    in_4 => mult3_p_net,
    in_5 => mult4_p_net,
    in_6 => mult5_p_net,
    in_7 => mult6_p_net,
    in_8 => mult7_p_net,
    in_9 => mult8_p_net,
    in_10 => mult9_p_net,
    in_11 => mult10_p_net,
    in_12 => mult11_p_net,
    in_13 => mult12_p_net,
    in_14 => mult13_p_net,
    in_15 => mult14_p_net,
    in_16 => mult15_p_net,
    out_1 => slice0_y_net_x1,
    out_2 => slice1_y_net_x1,
    out_3 => slice2_y_net_x1,
    out_4 => slice3_y_net_x1,
    out_5 => slice4_y_net_x1,
    out_6 => slice5_y_net_x1,
    out_7 => slice6_y_net_x1,
    out_8 => slice7_y_net_x1,
    out_9 => slice8_y_net_x1,
    out_10 => slice9_y_net_x1,
    out_11 => slice10_y_net_x1,
    out_12 => slice11_y_net_x1,
    out_13 => slice12_y_net_x1,
    out_14 => slice13_y_net_x1,
    out_15 => slice14_y_net_x1,
    out_16 => slice15_y_net_x1
  );
  vector_slice1 : entity xil_defaultlib.psb3_0_vector_slice1_x1 
  port map (
    in_1 => reinterpret0_output_port_net,
    in_2 => reinterpret1_output_port_net,
    in_3 => reinterpret2_output_port_net,
    in_4 => reinterpret3_output_port_net,
    in_5 => reinterpret4_output_port_net,
    in_6 => reinterpret5_output_port_net,
    in_7 => reinterpret6_output_port_net,
    in_8 => reinterpret7_output_port_net,
    in_9 => reinterpret8_output_port_net,
    in_10 => reinterpret9_output_port_net,
    in_11 => reinterpret10_output_port_net,
    in_12 => reinterpret11_output_port_net,
    in_13 => reinterpret12_output_port_net,
    in_14 => reinterpret13_output_port_net,
    in_15 => reinterpret14_output_port_net,
    in_16 => reinterpret15_output_port_net,
    out_1 => slice0_y_net_x0,
    out_2 => slice1_y_net_x0,
    out_3 => slice2_y_net_x0,
    out_4 => slice3_y_net_x0,
    out_5 => slice4_y_net_x0,
    out_6 => slice5_y_net_x0,
    out_7 => slice6_y_net_x0,
    out_8 => slice7_y_net_x0,
    out_9 => slice8_y_net_x0,
    out_10 => slice9_y_net_x0,
    out_11 => slice10_y_net_x0,
    out_12 => slice11_y_net_x0,
    out_13 => slice12_y_net_x0,
    out_14 => slice13_y_net_x0,
    out_15 => slice14_y_net_x0,
    out_16 => slice15_y_net_x0
  );
  vector_slice2 : entity xil_defaultlib.psb3_0_vector_slice2_x1 
  port map (
    in_1 => addsub0_s_net,
    in_2 => addsub1_s_net,
    in_3 => addsub2_s_net,
    in_4 => addsub3_s_net,
    in_5 => addsub4_s_net,
    in_6 => addsub5_s_net,
    in_7 => addsub6_s_net,
    in_8 => addsub7_s_net,
    in_9 => addsub8_s_net,
    in_10 => addsub9_s_net,
    in_11 => addsub10_s_net,
    in_12 => addsub11_s_net,
    in_13 => addsub12_s_net,
    in_14 => addsub13_s_net,
    in_15 => addsub14_s_net,
    in_16 => addsub15_s_net,
    out_1 => slice0_y_net,
    out_2 => slice1_y_net,
    out_3 => slice2_y_net,
    out_4 => slice3_y_net,
    out_5 => slice4_y_net,
    out_6 => slice5_y_net,
    out_7 => slice6_y_net,
    out_8 => slice7_y_net,
    out_9 => slice8_y_net,
    out_10 => slice9_y_net,
    out_11 => slice10_y_net,
    out_12 => slice11_y_net,
    out_13 => slice12_y_net,
    out_14 => slice13_y_net,
    out_15 => slice14_y_net,
    out_16 => slice15_y_net
  );
  vector_to_scalar : entity xil_defaultlib.psb3_0_vector_to_scalar_x1 
  port map (
    i_1 => delay0_q_net_x0,
    i_2 => delay1_q_net_x0,
    i_3 => delay2_q_net_x0,
    i_4 => delay3_q_net_x0,
    i_5 => delay4_q_net_x0,
    i_6 => delay5_q_net_x0,
    i_7 => delay6_q_net_x0,
    i_8 => delay7_q_net_x0,
    i_9 => delay8_q_net_x0,
    i_10 => delay9_q_net_x0,
    i_11 => delay10_q_net_x0,
    i_12 => delay11_q_net_x0,
    i_13 => delay12_q_net_x0,
    i_14 => delay13_q_net_x0,
    i_15 => delay14_q_net_x0,
    i_16 => delay15_q_net_x0,
    o => concat1_y_net_x1
  );
  vector_to_scalar1 : entity xil_defaultlib.psb3_0_vector_to_scalar1_x1 
  port map (
    i_1 => delay0_q_net,
    i_2 => delay1_q_net,
    i_3 => delay2_q_net,
    i_4 => delay3_q_net,
    i_5 => delay4_q_net,
    i_6 => delay5_q_net,
    i_7 => delay6_q_net,
    i_8 => delay7_q_net,
    i_9 => delay8_q_net,
    i_10 => delay9_q_net,
    i_11 => delay10_q_net,
    i_12 => delay11_q_net,
    i_13 => delay12_q_net,
    i_14 => delay13_q_net,
    i_15 => delay14_q_net,
    i_16 => delay15_q_net,
    o => concat1_y_net_x0
  );
  vector_to_scalar2 : entity xil_defaultlib.psb3_0_vector_to_scalar2 
  port map (
    i_1 => slice0_y_net,
    i_2 => slice1_y_net,
    i_3 => slice2_y_net,
    i_4 => slice3_y_net,
    i_5 => slice4_y_net,
    i_6 => slice5_y_net,
    i_7 => slice6_y_net,
    i_8 => slice7_y_net,
    i_9 => slice8_y_net,
    i_10 => slice9_y_net,
    i_11 => slice10_y_net,
    i_12 => slice11_y_net,
    i_13 => slice12_y_net,
    i_14 => slice13_y_net,
    i_15 => slice14_y_net,
    i_16 => slice15_y_net,
    o => concat1_y_net
  );
  constant17 : entity xil_defaultlib.sysgen_constant_71e89d757c 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant17_op_net
  );
  convert : entity xil_defaultlib.psb3_0_xlconvert 
  generic map (
    bool_conversion => 1,
    din_arith => 1,
    din_bin_pt => 0,
    din_width => 1,
    dout_arith => 1,
    dout_bin_pt => 0,
    dout_width => 1,
    latency => 1,
    overflow => xlWrap,
    quantization => xlTruncate
  )
  port map (
    clr => '0',
    en => "1",
    din => expression_dout_net,
    clk => clk_net,
    ce => ce_net,
    dout => convert_dout_net
  );
  expression : entity xil_defaultlib.sysgen_expr_7c83532765 
  port map (
    clr => '0',
    a => concat1_y_net_x1,
    b => concat1_y_net_x0,
    s => concat1_y_net,
    clk => clk_net,
    ce => ce_net,
    dout => expression_dout_net
  );
  register_x0 : entity xil_defaultlib.psb3_0_xlregister 
  generic map (
    d_width => 1,
    init_value => b"0"
  )
  port map (
    d => constant17_op_net,
    rst => gin_tl_reset_net,
    en => convert_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => register_q_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Overflow Detector add_im_4/Vector Delay
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_delay_x2 is
  port (
    d_1 : in std_logic_vector( 1-1 downto 0 );
    d_2 : in std_logic_vector( 1-1 downto 0 );
    d_3 : in std_logic_vector( 1-1 downto 0 );
    d_4 : in std_logic_vector( 1-1 downto 0 );
    d_5 : in std_logic_vector( 1-1 downto 0 );
    d_6 : in std_logic_vector( 1-1 downto 0 );
    d_7 : in std_logic_vector( 1-1 downto 0 );
    d_8 : in std_logic_vector( 1-1 downto 0 );
    d_9 : in std_logic_vector( 1-1 downto 0 );
    d_10 : in std_logic_vector( 1-1 downto 0 );
    d_11 : in std_logic_vector( 1-1 downto 0 );
    d_12 : in std_logic_vector( 1-1 downto 0 );
    d_13 : in std_logic_vector( 1-1 downto 0 );
    d_14 : in std_logic_vector( 1-1 downto 0 );
    d_15 : in std_logic_vector( 1-1 downto 0 );
    d_16 : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    q_1 : out std_logic_vector( 1-1 downto 0 );
    q_2 : out std_logic_vector( 1-1 downto 0 );
    q_3 : out std_logic_vector( 1-1 downto 0 );
    q_4 : out std_logic_vector( 1-1 downto 0 );
    q_5 : out std_logic_vector( 1-1 downto 0 );
    q_6 : out std_logic_vector( 1-1 downto 0 );
    q_7 : out std_logic_vector( 1-1 downto 0 );
    q_8 : out std_logic_vector( 1-1 downto 0 );
    q_9 : out std_logic_vector( 1-1 downto 0 );
    q_10 : out std_logic_vector( 1-1 downto 0 );
    q_11 : out std_logic_vector( 1-1 downto 0 );
    q_12 : out std_logic_vector( 1-1 downto 0 );
    q_13 : out std_logic_vector( 1-1 downto 0 );
    q_14 : out std_logic_vector( 1-1 downto 0 );
    q_15 : out std_logic_vector( 1-1 downto 0 );
    q_16 : out std_logic_vector( 1-1 downto 0 )
  );
end psb3_0_vector_delay_x2;
architecture structural of psb3_0_vector_delay_x2 is 
  signal delay4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay7_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay0_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay9_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay10_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay12_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay13_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay11_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal slice11_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay14_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal slice6_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay15_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 1-1 downto 0 );
begin
  q_1 <= delay0_q_net;
  q_2 <= delay1_q_net;
  q_3 <= delay2_q_net;
  q_4 <= delay3_q_net;
  q_5 <= delay4_q_net;
  q_6 <= delay5_q_net;
  q_7 <= delay6_q_net;
  q_8 <= delay7_q_net;
  q_9 <= delay8_q_net;
  q_10 <= delay9_q_net;
  q_11 <= delay10_q_net;
  q_12 <= delay11_q_net;
  q_13 <= delay12_q_net;
  q_14 <= delay13_q_net;
  q_15 <= delay14_q_net;
  q_16 <= delay15_q_net;
  slice0_y_net <= d_1;
  slice1_y_net <= d_2;
  slice2_y_net <= d_3;
  slice3_y_net <= d_4;
  slice4_y_net <= d_5;
  slice5_y_net <= d_6;
  slice6_y_net <= d_7;
  slice7_y_net <= d_8;
  slice8_y_net <= d_9;
  slice9_y_net <= d_10;
  slice10_y_net <= d_11;
  slice11_y_net <= d_12;
  slice12_y_net <= d_13;
  slice13_y_net <= d_14;
  slice14_y_net <= d_15;
  slice15_y_net <= d_16;
  clk_net <= clk_1;
  ce_net <= ce_1;
  delay0 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice0_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay0_q_net
  );
  delay1 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice2_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay3 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice3_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  delay4 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice4_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net
  );
  delay5 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice5_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  delay6 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice6_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay6_q_net
  );
  delay7 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice7_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay7_q_net
  );
  delay8 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice8_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay8_q_net
  );
  delay9 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice9_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay9_q_net
  );
  delay10 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice10_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay10_q_net
  );
  delay11 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice11_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay11_q_net
  );
  delay12 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice12_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay12_q_net
  );
  delay13 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice13_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay13_q_net
  );
  delay14 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice14_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay14_q_net
  );
  delay15 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice15_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay15_q_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Overflow Detector add_im_4/Vector Delay1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_delay1_x2 is
  port (
    d_1 : in std_logic_vector( 1-1 downto 0 );
    d_2 : in std_logic_vector( 1-1 downto 0 );
    d_3 : in std_logic_vector( 1-1 downto 0 );
    d_4 : in std_logic_vector( 1-1 downto 0 );
    d_5 : in std_logic_vector( 1-1 downto 0 );
    d_6 : in std_logic_vector( 1-1 downto 0 );
    d_7 : in std_logic_vector( 1-1 downto 0 );
    d_8 : in std_logic_vector( 1-1 downto 0 );
    d_9 : in std_logic_vector( 1-1 downto 0 );
    d_10 : in std_logic_vector( 1-1 downto 0 );
    d_11 : in std_logic_vector( 1-1 downto 0 );
    d_12 : in std_logic_vector( 1-1 downto 0 );
    d_13 : in std_logic_vector( 1-1 downto 0 );
    d_14 : in std_logic_vector( 1-1 downto 0 );
    d_15 : in std_logic_vector( 1-1 downto 0 );
    d_16 : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    q_1 : out std_logic_vector( 1-1 downto 0 );
    q_2 : out std_logic_vector( 1-1 downto 0 );
    q_3 : out std_logic_vector( 1-1 downto 0 );
    q_4 : out std_logic_vector( 1-1 downto 0 );
    q_5 : out std_logic_vector( 1-1 downto 0 );
    q_6 : out std_logic_vector( 1-1 downto 0 );
    q_7 : out std_logic_vector( 1-1 downto 0 );
    q_8 : out std_logic_vector( 1-1 downto 0 );
    q_9 : out std_logic_vector( 1-1 downto 0 );
    q_10 : out std_logic_vector( 1-1 downto 0 );
    q_11 : out std_logic_vector( 1-1 downto 0 );
    q_12 : out std_logic_vector( 1-1 downto 0 );
    q_13 : out std_logic_vector( 1-1 downto 0 );
    q_14 : out std_logic_vector( 1-1 downto 0 );
    q_15 : out std_logic_vector( 1-1 downto 0 );
    q_16 : out std_logic_vector( 1-1 downto 0 )
  );
end psb3_0_vector_delay1_x2;
architecture structural of psb3_0_vector_delay1_x2 is 
  signal delay0_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay13_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay12_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay7_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay9_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay14_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay15_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay10_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay11_q_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal slice13_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
begin
  q_1 <= delay0_q_net;
  q_2 <= delay1_q_net;
  q_3 <= delay2_q_net;
  q_4 <= delay3_q_net;
  q_5 <= delay4_q_net;
  q_6 <= delay5_q_net;
  q_7 <= delay6_q_net;
  q_8 <= delay7_q_net;
  q_9 <= delay8_q_net;
  q_10 <= delay9_q_net;
  q_11 <= delay10_q_net;
  q_12 <= delay11_q_net;
  q_13 <= delay12_q_net;
  q_14 <= delay13_q_net;
  q_15 <= delay14_q_net;
  q_16 <= delay15_q_net;
  slice0_y_net <= d_1;
  slice1_y_net <= d_2;
  slice2_y_net <= d_3;
  slice3_y_net <= d_4;
  slice4_y_net <= d_5;
  slice5_y_net <= d_6;
  slice6_y_net <= d_7;
  slice7_y_net <= d_8;
  slice8_y_net <= d_9;
  slice9_y_net <= d_10;
  slice10_y_net <= d_11;
  slice11_y_net <= d_12;
  slice12_y_net <= d_13;
  slice13_y_net <= d_14;
  slice14_y_net <= d_15;
  slice15_y_net <= d_16;
  clk_net <= clk_1;
  ce_net <= ce_1;
  delay0 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice0_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay0_q_net
  );
  delay1 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice2_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay3 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice3_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  delay4 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice4_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net
  );
  delay5 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice5_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  delay6 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice6_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay6_q_net
  );
  delay7 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice7_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay7_q_net
  );
  delay8 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice8_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay8_q_net
  );
  delay9 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice9_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay9_q_net
  );
  delay10 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice10_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay10_q_net
  );
  delay11 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice11_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay11_q_net
  );
  delay12 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice12_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay12_q_net
  );
  delay13 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice13_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay13_q_net
  );
  delay14 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice14_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay14_q_net
  );
  delay15 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice15_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay15_q_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Overflow Detector add_im_4/Vector Slice
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_slice_x2 is
  port (
    in_1 : in std_logic_vector( 16-1 downto 0 );
    in_2 : in std_logic_vector( 16-1 downto 0 );
    in_3 : in std_logic_vector( 16-1 downto 0 );
    in_4 : in std_logic_vector( 16-1 downto 0 );
    in_5 : in std_logic_vector( 16-1 downto 0 );
    in_6 : in std_logic_vector( 16-1 downto 0 );
    in_7 : in std_logic_vector( 16-1 downto 0 );
    in_8 : in std_logic_vector( 16-1 downto 0 );
    in_9 : in std_logic_vector( 16-1 downto 0 );
    in_10 : in std_logic_vector( 16-1 downto 0 );
    in_11 : in std_logic_vector( 16-1 downto 0 );
    in_12 : in std_logic_vector( 16-1 downto 0 );
    in_13 : in std_logic_vector( 16-1 downto 0 );
    in_14 : in std_logic_vector( 16-1 downto 0 );
    in_15 : in std_logic_vector( 16-1 downto 0 );
    in_16 : in std_logic_vector( 16-1 downto 0 );
    out_1 : out std_logic_vector( 1-1 downto 0 );
    out_2 : out std_logic_vector( 1-1 downto 0 );
    out_3 : out std_logic_vector( 1-1 downto 0 );
    out_4 : out std_logic_vector( 1-1 downto 0 );
    out_5 : out std_logic_vector( 1-1 downto 0 );
    out_6 : out std_logic_vector( 1-1 downto 0 );
    out_7 : out std_logic_vector( 1-1 downto 0 );
    out_8 : out std_logic_vector( 1-1 downto 0 );
    out_9 : out std_logic_vector( 1-1 downto 0 );
    out_10 : out std_logic_vector( 1-1 downto 0 );
    out_11 : out std_logic_vector( 1-1 downto 0 );
    out_12 : out std_logic_vector( 1-1 downto 0 );
    out_13 : out std_logic_vector( 1-1 downto 0 );
    out_14 : out std_logic_vector( 1-1 downto 0 );
    out_15 : out std_logic_vector( 1-1 downto 0 );
    out_16 : out std_logic_vector( 1-1 downto 0 )
  );
end psb3_0_vector_slice_x2;
architecture structural of psb3_0_vector_slice_x2 is 
  signal slice6_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 1-1 downto 0 );
  signal mult10_p_net : std_logic_vector( 16-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 1-1 downto 0 );
  signal mult2_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult1_p_net : std_logic_vector( 16-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 1-1 downto 0 );
  signal mult4_p_net : std_logic_vector( 16-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 1-1 downto 0 );
  signal mult6_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult13_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult0_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult12_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult15_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult11_p_net : std_logic_vector( 16-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 1-1 downto 0 );
  signal mult3_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult7_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult9_p_net : std_logic_vector( 16-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 1-1 downto 0 );
  signal mult14_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult5_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult8_p_net : std_logic_vector( 16-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 1-1 downto 0 );
begin
  out_1 <= slice0_y_net;
  out_2 <= slice1_y_net;
  out_3 <= slice2_y_net;
  out_4 <= slice3_y_net;
  out_5 <= slice4_y_net;
  out_6 <= slice5_y_net;
  out_7 <= slice6_y_net;
  out_8 <= slice7_y_net;
  out_9 <= slice8_y_net;
  out_10 <= slice9_y_net;
  out_11 <= slice10_y_net;
  out_12 <= slice11_y_net;
  out_13 <= slice12_y_net;
  out_14 <= slice13_y_net;
  out_15 <= slice14_y_net;
  out_16 <= slice15_y_net;
  mult0_p_net <= in_1;
  mult1_p_net <= in_2;
  mult2_p_net <= in_3;
  mult3_p_net <= in_4;
  mult4_p_net <= in_5;
  mult5_p_net <= in_6;
  mult6_p_net <= in_7;
  mult7_p_net <= in_8;
  mult8_p_net <= in_9;
  mult9_p_net <= in_10;
  mult10_p_net <= in_11;
  mult11_p_net <= in_12;
  mult12_p_net <= in_13;
  mult13_p_net <= in_14;
  mult14_p_net <= in_15;
  mult15_p_net <= in_16;
  slice0 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult0_p_net,
    y => slice0_y_net
  );
  slice1 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult1_p_net,
    y => slice1_y_net
  );
  slice2 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult2_p_net,
    y => slice2_y_net
  );
  slice3 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult3_p_net,
    y => slice3_y_net
  );
  slice4 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult4_p_net,
    y => slice4_y_net
  );
  slice5 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult5_p_net,
    y => slice5_y_net
  );
  slice6 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult6_p_net,
    y => slice6_y_net
  );
  slice7 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult7_p_net,
    y => slice7_y_net
  );
  slice8 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult8_p_net,
    y => slice8_y_net
  );
  slice9 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult9_p_net,
    y => slice9_y_net
  );
  slice10 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult10_p_net,
    y => slice10_y_net
  );
  slice11 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult11_p_net,
    y => slice11_y_net
  );
  slice12 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult12_p_net,
    y => slice12_y_net
  );
  slice13 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult13_p_net,
    y => slice13_y_net
  );
  slice14 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult14_p_net,
    y => slice14_y_net
  );
  slice15 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult15_p_net,
    y => slice15_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Overflow Detector add_im_4/Vector Slice1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_slice1_x2 is
  port (
    in_1 : in std_logic_vector( 16-1 downto 0 );
    in_2 : in std_logic_vector( 16-1 downto 0 );
    in_3 : in std_logic_vector( 16-1 downto 0 );
    in_4 : in std_logic_vector( 16-1 downto 0 );
    in_5 : in std_logic_vector( 16-1 downto 0 );
    in_6 : in std_logic_vector( 16-1 downto 0 );
    in_7 : in std_logic_vector( 16-1 downto 0 );
    in_8 : in std_logic_vector( 16-1 downto 0 );
    in_9 : in std_logic_vector( 16-1 downto 0 );
    in_10 : in std_logic_vector( 16-1 downto 0 );
    in_11 : in std_logic_vector( 16-1 downto 0 );
    in_12 : in std_logic_vector( 16-1 downto 0 );
    in_13 : in std_logic_vector( 16-1 downto 0 );
    in_14 : in std_logic_vector( 16-1 downto 0 );
    in_15 : in std_logic_vector( 16-1 downto 0 );
    in_16 : in std_logic_vector( 16-1 downto 0 );
    out_1 : out std_logic_vector( 1-1 downto 0 );
    out_2 : out std_logic_vector( 1-1 downto 0 );
    out_3 : out std_logic_vector( 1-1 downto 0 );
    out_4 : out std_logic_vector( 1-1 downto 0 );
    out_5 : out std_logic_vector( 1-1 downto 0 );
    out_6 : out std_logic_vector( 1-1 downto 0 );
    out_7 : out std_logic_vector( 1-1 downto 0 );
    out_8 : out std_logic_vector( 1-1 downto 0 );
    out_9 : out std_logic_vector( 1-1 downto 0 );
    out_10 : out std_logic_vector( 1-1 downto 0 );
    out_11 : out std_logic_vector( 1-1 downto 0 );
    out_12 : out std_logic_vector( 1-1 downto 0 );
    out_13 : out std_logic_vector( 1-1 downto 0 );
    out_14 : out std_logic_vector( 1-1 downto 0 );
    out_15 : out std_logic_vector( 1-1 downto 0 );
    out_16 : out std_logic_vector( 1-1 downto 0 )
  );
end psb3_0_vector_slice1_x2;
architecture structural of psb3_0_vector_slice1_x2 is 
  signal slice15_y_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
begin
  out_1 <= slice0_y_net;
  out_2 <= slice1_y_net;
  out_3 <= slice2_y_net;
  out_4 <= slice3_y_net;
  out_5 <= slice4_y_net;
  out_6 <= slice5_y_net;
  out_7 <= slice6_y_net;
  out_8 <= slice7_y_net;
  out_9 <= slice8_y_net;
  out_10 <= slice9_y_net;
  out_11 <= slice10_y_net;
  out_12 <= slice11_y_net;
  out_13 <= slice12_y_net;
  out_14 <= slice13_y_net;
  out_15 <= slice14_y_net;
  out_16 <= slice15_y_net;
  reinterpret0_output_port_net <= in_1;
  reinterpret1_output_port_net <= in_2;
  reinterpret2_output_port_net <= in_3;
  reinterpret3_output_port_net <= in_4;
  reinterpret4_output_port_net <= in_5;
  reinterpret5_output_port_net <= in_6;
  reinterpret6_output_port_net <= in_7;
  reinterpret7_output_port_net <= in_8;
  reinterpret8_output_port_net <= in_9;
  reinterpret9_output_port_net <= in_10;
  reinterpret10_output_port_net <= in_11;
  reinterpret11_output_port_net <= in_12;
  reinterpret12_output_port_net <= in_13;
  reinterpret13_output_port_net <= in_14;
  reinterpret14_output_port_net <= in_15;
  reinterpret15_output_port_net <= in_16;
  slice0 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret0_output_port_net,
    y => slice0_y_net
  );
  slice1 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret1_output_port_net,
    y => slice1_y_net
  );
  slice2 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret2_output_port_net,
    y => slice2_y_net
  );
  slice3 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret3_output_port_net,
    y => slice3_y_net
  );
  slice4 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret4_output_port_net,
    y => slice4_y_net
  );
  slice5 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret5_output_port_net,
    y => slice5_y_net
  );
  slice6 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret6_output_port_net,
    y => slice6_y_net
  );
  slice7 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret7_output_port_net,
    y => slice7_y_net
  );
  slice8 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret8_output_port_net,
    y => slice8_y_net
  );
  slice9 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret9_output_port_net,
    y => slice9_y_net
  );
  slice10 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret10_output_port_net,
    y => slice10_y_net
  );
  slice11 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret11_output_port_net,
    y => slice11_y_net
  );
  slice12 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret12_output_port_net,
    y => slice12_y_net
  );
  slice13 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret13_output_port_net,
    y => slice13_y_net
  );
  slice14 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret14_output_port_net,
    y => slice14_y_net
  );
  slice15 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret15_output_port_net,
    y => slice15_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Overflow Detector add_im_4/Vector Slice2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_slice2_x2 is
  port (
    in_1 : in std_logic_vector( 16-1 downto 0 );
    in_2 : in std_logic_vector( 16-1 downto 0 );
    in_3 : in std_logic_vector( 16-1 downto 0 );
    in_4 : in std_logic_vector( 16-1 downto 0 );
    in_5 : in std_logic_vector( 16-1 downto 0 );
    in_6 : in std_logic_vector( 16-1 downto 0 );
    in_7 : in std_logic_vector( 16-1 downto 0 );
    in_8 : in std_logic_vector( 16-1 downto 0 );
    in_9 : in std_logic_vector( 16-1 downto 0 );
    in_10 : in std_logic_vector( 16-1 downto 0 );
    in_11 : in std_logic_vector( 16-1 downto 0 );
    in_12 : in std_logic_vector( 16-1 downto 0 );
    in_13 : in std_logic_vector( 16-1 downto 0 );
    in_14 : in std_logic_vector( 16-1 downto 0 );
    in_15 : in std_logic_vector( 16-1 downto 0 );
    in_16 : in std_logic_vector( 16-1 downto 0 );
    out_1 : out std_logic_vector( 1-1 downto 0 );
    out_2 : out std_logic_vector( 1-1 downto 0 );
    out_3 : out std_logic_vector( 1-1 downto 0 );
    out_4 : out std_logic_vector( 1-1 downto 0 );
    out_5 : out std_logic_vector( 1-1 downto 0 );
    out_6 : out std_logic_vector( 1-1 downto 0 );
    out_7 : out std_logic_vector( 1-1 downto 0 );
    out_8 : out std_logic_vector( 1-1 downto 0 );
    out_9 : out std_logic_vector( 1-1 downto 0 );
    out_10 : out std_logic_vector( 1-1 downto 0 );
    out_11 : out std_logic_vector( 1-1 downto 0 );
    out_12 : out std_logic_vector( 1-1 downto 0 );
    out_13 : out std_logic_vector( 1-1 downto 0 );
    out_14 : out std_logic_vector( 1-1 downto 0 );
    out_15 : out std_logic_vector( 1-1 downto 0 );
    out_16 : out std_logic_vector( 1-1 downto 0 )
  );
end psb3_0_vector_slice2_x2;
architecture structural of psb3_0_vector_slice2_x2 is 
  signal slice1_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 1-1 downto 0 );
  signal addsub11_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub7_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub8_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub9_s_net : std_logic_vector( 16-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 1-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub0_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub6_s_net : std_logic_vector( 16-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 1-1 downto 0 );
  signal addsub12_s_net : std_logic_vector( 16-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 1-1 downto 0 );
  signal addsub15_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub13_s_net : std_logic_vector( 16-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 1-1 downto 0 );
  signal addsub3_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub5_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub10_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub14_s_net : std_logic_vector( 16-1 downto 0 );
begin
  out_1 <= slice0_y_net;
  out_2 <= slice1_y_net;
  out_3 <= slice2_y_net;
  out_4 <= slice3_y_net;
  out_5 <= slice4_y_net;
  out_6 <= slice5_y_net;
  out_7 <= slice6_y_net;
  out_8 <= slice7_y_net;
  out_9 <= slice8_y_net;
  out_10 <= slice9_y_net;
  out_11 <= slice10_y_net;
  out_12 <= slice11_y_net;
  out_13 <= slice12_y_net;
  out_14 <= slice13_y_net;
  out_15 <= slice14_y_net;
  out_16 <= slice15_y_net;
  addsub0_s_net <= in_1;
  addsub1_s_net <= in_2;
  addsub2_s_net <= in_3;
  addsub3_s_net <= in_4;
  addsub4_s_net <= in_5;
  addsub5_s_net <= in_6;
  addsub6_s_net <= in_7;
  addsub7_s_net <= in_8;
  addsub8_s_net <= in_9;
  addsub9_s_net <= in_10;
  addsub10_s_net <= in_11;
  addsub11_s_net <= in_12;
  addsub12_s_net <= in_13;
  addsub13_s_net <= in_14;
  addsub14_s_net <= in_15;
  addsub15_s_net <= in_16;
  slice0 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub0_s_net,
    y => slice0_y_net
  );
  slice1 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub1_s_net,
    y => slice1_y_net
  );
  slice2 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub2_s_net,
    y => slice2_y_net
  );
  slice3 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub3_s_net,
    y => slice3_y_net
  );
  slice4 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub4_s_net,
    y => slice4_y_net
  );
  slice5 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub5_s_net,
    y => slice5_y_net
  );
  slice6 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub6_s_net,
    y => slice6_y_net
  );
  slice7 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub7_s_net,
    y => slice7_y_net
  );
  slice8 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub8_s_net,
    y => slice8_y_net
  );
  slice9 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub9_s_net,
    y => slice9_y_net
  );
  slice10 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub10_s_net,
    y => slice10_y_net
  );
  slice11 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub11_s_net,
    y => slice11_y_net
  );
  slice12 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub12_s_net,
    y => slice12_y_net
  );
  slice13 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub13_s_net,
    y => slice13_y_net
  );
  slice14 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub14_s_net,
    y => slice14_y_net
  );
  slice15 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub15_s_net,
    y => slice15_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Overflow Detector add_im_4/Vector to Scalar
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_to_scalar_x2 is
  port (
    i_1 : in std_logic_vector( 1-1 downto 0 );
    i_2 : in std_logic_vector( 1-1 downto 0 );
    i_3 : in std_logic_vector( 1-1 downto 0 );
    i_4 : in std_logic_vector( 1-1 downto 0 );
    i_5 : in std_logic_vector( 1-1 downto 0 );
    i_6 : in std_logic_vector( 1-1 downto 0 );
    i_7 : in std_logic_vector( 1-1 downto 0 );
    i_8 : in std_logic_vector( 1-1 downto 0 );
    i_9 : in std_logic_vector( 1-1 downto 0 );
    i_10 : in std_logic_vector( 1-1 downto 0 );
    i_11 : in std_logic_vector( 1-1 downto 0 );
    i_12 : in std_logic_vector( 1-1 downto 0 );
    i_13 : in std_logic_vector( 1-1 downto 0 );
    i_14 : in std_logic_vector( 1-1 downto 0 );
    i_15 : in std_logic_vector( 1-1 downto 0 );
    i_16 : in std_logic_vector( 1-1 downto 0 );
    o : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_vector_to_scalar_x2;
architecture structural of psb3_0_vector_to_scalar_x2 is 
  signal delay5_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay11_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay9_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay12_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay13_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay14_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay15_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay10_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay7_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay0_q_net : std_logic_vector( 1-1 downto 0 );
  signal concat1_y_net : std_logic_vector( 16-1 downto 0 );
begin
  o <= concat1_y_net;
  delay0_q_net <= i_1;
  delay1_q_net <= i_2;
  delay2_q_net <= i_3;
  delay3_q_net <= i_4;
  delay4_q_net <= i_5;
  delay5_q_net <= i_6;
  delay6_q_net <= i_7;
  delay7_q_net <= i_8;
  delay8_q_net <= i_9;
  delay9_q_net <= i_10;
  delay10_q_net <= i_11;
  delay11_q_net <= i_12;
  delay12_q_net <= i_13;
  delay13_q_net <= i_14;
  delay14_q_net <= i_15;
  delay15_q_net <= i_16;
  concat1 : entity xil_defaultlib.sysgen_concat_d977c66e35 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => delay15_q_net,
    in1 => delay14_q_net,
    in2 => delay13_q_net,
    in3 => delay12_q_net,
    in4 => delay11_q_net,
    in5 => delay10_q_net,
    in6 => delay9_q_net,
    in7 => delay8_q_net,
    in8 => delay7_q_net,
    in9 => delay6_q_net,
    in10 => delay5_q_net,
    in11 => delay4_q_net,
    in12 => delay3_q_net,
    in13 => delay2_q_net,
    in14 => delay1_q_net,
    in15 => delay0_q_net,
    y => concat1_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Overflow Detector add_im_4/Vector to Scalar1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_to_scalar1_x2 is
  port (
    i_1 : in std_logic_vector( 1-1 downto 0 );
    i_2 : in std_logic_vector( 1-1 downto 0 );
    i_3 : in std_logic_vector( 1-1 downto 0 );
    i_4 : in std_logic_vector( 1-1 downto 0 );
    i_5 : in std_logic_vector( 1-1 downto 0 );
    i_6 : in std_logic_vector( 1-1 downto 0 );
    i_7 : in std_logic_vector( 1-1 downto 0 );
    i_8 : in std_logic_vector( 1-1 downto 0 );
    i_9 : in std_logic_vector( 1-1 downto 0 );
    i_10 : in std_logic_vector( 1-1 downto 0 );
    i_11 : in std_logic_vector( 1-1 downto 0 );
    i_12 : in std_logic_vector( 1-1 downto 0 );
    i_13 : in std_logic_vector( 1-1 downto 0 );
    i_14 : in std_logic_vector( 1-1 downto 0 );
    i_15 : in std_logic_vector( 1-1 downto 0 );
    i_16 : in std_logic_vector( 1-1 downto 0 );
    o : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_vector_to_scalar1_x2;
architecture structural of psb3_0_vector_to_scalar1_x2 is 
  signal delay14_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay7_q_net : std_logic_vector( 1-1 downto 0 );
  signal concat1_y_net : std_logic_vector( 16-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay13_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay10_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay15_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay12_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay0_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay9_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay11_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
begin
  o <= concat1_y_net;
  delay0_q_net <= i_1;
  delay1_q_net <= i_2;
  delay2_q_net <= i_3;
  delay3_q_net <= i_4;
  delay4_q_net <= i_5;
  delay5_q_net <= i_6;
  delay6_q_net <= i_7;
  delay7_q_net <= i_8;
  delay8_q_net <= i_9;
  delay9_q_net <= i_10;
  delay10_q_net <= i_11;
  delay11_q_net <= i_12;
  delay12_q_net <= i_13;
  delay13_q_net <= i_14;
  delay14_q_net <= i_15;
  delay15_q_net <= i_16;
  concat1 : entity xil_defaultlib.sysgen_concat_d977c66e35 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => delay15_q_net,
    in1 => delay14_q_net,
    in2 => delay13_q_net,
    in3 => delay12_q_net,
    in4 => delay11_q_net,
    in5 => delay10_q_net,
    in6 => delay9_q_net,
    in7 => delay8_q_net,
    in8 => delay7_q_net,
    in9 => delay6_q_net,
    in10 => delay5_q_net,
    in11 => delay4_q_net,
    in12 => delay3_q_net,
    in13 => delay2_q_net,
    in14 => delay1_q_net,
    in15 => delay0_q_net,
    y => concat1_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Overflow Detector add_im_4/Vector to Scalar2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_to_scalar2_x2 is
  port (
    i_1 : in std_logic_vector( 1-1 downto 0 );
    i_2 : in std_logic_vector( 1-1 downto 0 );
    i_3 : in std_logic_vector( 1-1 downto 0 );
    i_4 : in std_logic_vector( 1-1 downto 0 );
    i_5 : in std_logic_vector( 1-1 downto 0 );
    i_6 : in std_logic_vector( 1-1 downto 0 );
    i_7 : in std_logic_vector( 1-1 downto 0 );
    i_8 : in std_logic_vector( 1-1 downto 0 );
    i_9 : in std_logic_vector( 1-1 downto 0 );
    i_10 : in std_logic_vector( 1-1 downto 0 );
    i_11 : in std_logic_vector( 1-1 downto 0 );
    i_12 : in std_logic_vector( 1-1 downto 0 );
    i_13 : in std_logic_vector( 1-1 downto 0 );
    i_14 : in std_logic_vector( 1-1 downto 0 );
    i_15 : in std_logic_vector( 1-1 downto 0 );
    i_16 : in std_logic_vector( 1-1 downto 0 );
    o : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_vector_to_scalar2_x2;
architecture structural of psb3_0_vector_to_scalar2_x2 is 
  signal concat1_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 1-1 downto 0 );
begin
  o <= concat1_y_net;
  slice0_y_net <= i_1;
  slice1_y_net <= i_2;
  slice2_y_net <= i_3;
  slice3_y_net <= i_4;
  slice4_y_net <= i_5;
  slice5_y_net <= i_6;
  slice6_y_net <= i_7;
  slice7_y_net <= i_8;
  slice8_y_net <= i_9;
  slice9_y_net <= i_10;
  slice10_y_net <= i_11;
  slice11_y_net <= i_12;
  slice12_y_net <= i_13;
  slice13_y_net <= i_14;
  slice14_y_net <= i_15;
  slice15_y_net <= i_16;
  concat1 : entity xil_defaultlib.sysgen_concat_d977c66e35 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => slice15_y_net,
    in1 => slice14_y_net,
    in2 => slice13_y_net,
    in3 => slice12_y_net,
    in4 => slice11_y_net,
    in5 => slice10_y_net,
    in6 => slice9_y_net,
    in7 => slice8_y_net,
    in8 => slice7_y_net,
    in9 => slice6_y_net,
    in10 => slice5_y_net,
    in11 => slice4_y_net,
    in12 => slice3_y_net,
    in13 => slice2_y_net,
    in14 => slice1_y_net,
    in15 => slice0_y_net,
    y => concat1_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Overflow Detector add_im_4
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_overflow_detector_add_im_4 is
  port (
    rst : in std_logic_vector( 1-1 downto 0 );
    a_1 : in std_logic_vector( 16-1 downto 0 );
    b_1 : in std_logic_vector( 16-1 downto 0 );
    s_1 : in std_logic_vector( 16-1 downto 0 );
    a_2 : in std_logic_vector( 16-1 downto 0 );
    a_3 : in std_logic_vector( 16-1 downto 0 );
    a_4 : in std_logic_vector( 16-1 downto 0 );
    a_5 : in std_logic_vector( 16-1 downto 0 );
    a_6 : in std_logic_vector( 16-1 downto 0 );
    a_7 : in std_logic_vector( 16-1 downto 0 );
    a_8 : in std_logic_vector( 16-1 downto 0 );
    a_9 : in std_logic_vector( 16-1 downto 0 );
    a_10 : in std_logic_vector( 16-1 downto 0 );
    a_11 : in std_logic_vector( 16-1 downto 0 );
    a_12 : in std_logic_vector( 16-1 downto 0 );
    a_13 : in std_logic_vector( 16-1 downto 0 );
    a_14 : in std_logic_vector( 16-1 downto 0 );
    a_15 : in std_logic_vector( 16-1 downto 0 );
    a_16 : in std_logic_vector( 16-1 downto 0 );
    b_2 : in std_logic_vector( 16-1 downto 0 );
    b_3 : in std_logic_vector( 16-1 downto 0 );
    b_4 : in std_logic_vector( 16-1 downto 0 );
    b_5 : in std_logic_vector( 16-1 downto 0 );
    b_6 : in std_logic_vector( 16-1 downto 0 );
    b_7 : in std_logic_vector( 16-1 downto 0 );
    b_8 : in std_logic_vector( 16-1 downto 0 );
    b_9 : in std_logic_vector( 16-1 downto 0 );
    b_10 : in std_logic_vector( 16-1 downto 0 );
    b_11 : in std_logic_vector( 16-1 downto 0 );
    b_12 : in std_logic_vector( 16-1 downto 0 );
    b_13 : in std_logic_vector( 16-1 downto 0 );
    b_14 : in std_logic_vector( 16-1 downto 0 );
    b_15 : in std_logic_vector( 16-1 downto 0 );
    b_16 : in std_logic_vector( 16-1 downto 0 );
    s_2 : in std_logic_vector( 16-1 downto 0 );
    s_3 : in std_logic_vector( 16-1 downto 0 );
    s_4 : in std_logic_vector( 16-1 downto 0 );
    s_5 : in std_logic_vector( 16-1 downto 0 );
    s_6 : in std_logic_vector( 16-1 downto 0 );
    s_7 : in std_logic_vector( 16-1 downto 0 );
    s_8 : in std_logic_vector( 16-1 downto 0 );
    s_9 : in std_logic_vector( 16-1 downto 0 );
    s_10 : in std_logic_vector( 16-1 downto 0 );
    s_11 : in std_logic_vector( 16-1 downto 0 );
    s_12 : in std_logic_vector( 16-1 downto 0 );
    s_13 : in std_logic_vector( 16-1 downto 0 );
    s_14 : in std_logic_vector( 16-1 downto 0 );
    s_15 : in std_logic_vector( 16-1 downto 0 );
    s_16 : in std_logic_vector( 16-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    ov : out std_logic_vector( 1-1 downto 0 )
  );
end psb3_0_overflow_detector_add_im_4;
architecture structural of psb3_0_overflow_detector_add_im_4 is 
  signal addsub14_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 16-1 downto 0 );
  signal delay10_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay13_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal addsub11_s_net : std_logic_vector( 16-1 downto 0 );
  signal delay6_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice1_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal addsub8_s_net : std_logic_vector( 16-1 downto 0 );
  signal delay4_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay12_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice7_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal addsub15_s_net : std_logic_vector( 16-1 downto 0 );
  signal slice9_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 16-1 downto 0 );
  signal delay8_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice10_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal slice12_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal delay14_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay11_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice6_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal slice11_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal slice13_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal slice14_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal slice4_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal addsub5_s_net : std_logic_vector( 16-1 downto 0 );
  signal delay15_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice2_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal slice5_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal slice15_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal delay0_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal addsub13_s_net : std_logic_vector( 16-1 downto 0 );
  signal clk_net : std_logic;
  signal addsub3_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub7_s_net : std_logic_vector( 16-1 downto 0 );
  signal ce_net : std_logic;
  signal delay2_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal addsub9_s_net : std_logic_vector( 16-1 downto 0 );
  signal delay3_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal addsub6_s_net : std_logic_vector( 16-1 downto 0 );
  signal delay5_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay7_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay9_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal addsub12_s_net : std_logic_vector( 16-1 downto 0 );
  signal slice0_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal slice3_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal slice8_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal delay0_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal addsub10_s_net : std_logic_vector( 16-1 downto 0 );
  signal delay11_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay15_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice0_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice6_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice7_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice2_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice14_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay9_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice9_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice3_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice1_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay10_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 1-1 downto 0 );
  signal concat1_y_net_x1 : std_logic_vector( 16-1 downto 0 );
  signal constant17_op_net : std_logic_vector( 1-1 downto 0 );
  signal delay14_q_net : std_logic_vector( 1-1 downto 0 );
  signal concat1_y_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal delay12_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice13_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice4_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 1-1 downto 0 );
  signal concat1_y_net : std_logic_vector( 16-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice10_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice12_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay7_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay13_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice11_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice5_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal convert_dout_net : std_logic_vector( 1-1 downto 0 );
  signal expression_dout_net : std_logic_vector( 1-1 downto 0 );
  signal slice8_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice15_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal gin_tl_reset_net : std_logic_vector( 1-1 downto 0 );
  signal register_q_net : std_logic_vector( 1-1 downto 0 );
  signal mult0_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub0_s_net : std_logic_vector( 16-1 downto 0 );
  signal mult2_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult10_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult12_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mult14_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult13_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult6_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mult7_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult3_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mult8_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mult4_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mult11_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult1_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 16-1 downto 0 );
  signal mult5_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mult15_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult9_p_net : std_logic_vector( 16-1 downto 0 );
begin
  ov <= register_q_net;
  gin_tl_reset_net <= rst;
  mult0_p_net <= a_1;
  reinterpret0_output_port_net <= b_1;
  addsub0_s_net <= s_1;
  mult1_p_net <= a_2;
  mult2_p_net <= a_3;
  mult3_p_net <= a_4;
  mult4_p_net <= a_5;
  mult5_p_net <= a_6;
  mult6_p_net <= a_7;
  mult7_p_net <= a_8;
  mult8_p_net <= a_9;
  mult9_p_net <= a_10;
  mult10_p_net <= a_11;
  mult11_p_net <= a_12;
  mult12_p_net <= a_13;
  mult13_p_net <= a_14;
  mult14_p_net <= a_15;
  mult15_p_net <= a_16;
  reinterpret1_output_port_net <= b_2;
  reinterpret2_output_port_net <= b_3;
  reinterpret3_output_port_net <= b_4;
  reinterpret4_output_port_net <= b_5;
  reinterpret5_output_port_net <= b_6;
  reinterpret6_output_port_net <= b_7;
  reinterpret7_output_port_net <= b_8;
  reinterpret8_output_port_net <= b_9;
  reinterpret9_output_port_net <= b_10;
  reinterpret10_output_port_net <= b_11;
  reinterpret11_output_port_net <= b_12;
  reinterpret12_output_port_net <= b_13;
  reinterpret13_output_port_net <= b_14;
  reinterpret14_output_port_net <= b_15;
  reinterpret15_output_port_net <= b_16;
  addsub1_s_net <= s_2;
  addsub2_s_net <= s_3;
  addsub3_s_net <= s_4;
  addsub4_s_net <= s_5;
  addsub5_s_net <= s_6;
  addsub6_s_net <= s_7;
  addsub7_s_net <= s_8;
  addsub8_s_net <= s_9;
  addsub9_s_net <= s_10;
  addsub10_s_net <= s_11;
  addsub11_s_net <= s_12;
  addsub12_s_net <= s_13;
  addsub13_s_net <= s_14;
  addsub14_s_net <= s_15;
  addsub15_s_net <= s_16;
  clk_net <= clk_1;
  ce_net <= ce_1;
  vector_delay : entity xil_defaultlib.psb3_0_vector_delay_x2 
  port map (
    d_1 => slice0_y_net_x1,
    d_2 => slice1_y_net_x1,
    d_3 => slice2_y_net_x1,
    d_4 => slice3_y_net_x1,
    d_5 => slice4_y_net_x1,
    d_6 => slice5_y_net_x1,
    d_7 => slice6_y_net_x1,
    d_8 => slice7_y_net_x1,
    d_9 => slice8_y_net_x1,
    d_10 => slice9_y_net_x1,
    d_11 => slice10_y_net_x1,
    d_12 => slice11_y_net_x1,
    d_13 => slice12_y_net_x1,
    d_14 => slice13_y_net_x1,
    d_15 => slice14_y_net_x1,
    d_16 => slice15_y_net_x1,
    clk_1 => clk_net,
    ce_1 => ce_net,
    q_1 => delay0_q_net_x0,
    q_2 => delay1_q_net_x0,
    q_3 => delay2_q_net_x0,
    q_4 => delay3_q_net_x0,
    q_5 => delay4_q_net_x0,
    q_6 => delay5_q_net_x0,
    q_7 => delay6_q_net_x0,
    q_8 => delay7_q_net_x0,
    q_9 => delay8_q_net_x0,
    q_10 => delay9_q_net_x0,
    q_11 => delay10_q_net_x0,
    q_12 => delay11_q_net_x0,
    q_13 => delay12_q_net_x0,
    q_14 => delay13_q_net_x0,
    q_15 => delay14_q_net_x0,
    q_16 => delay15_q_net_x0
  );
  vector_delay1 : entity xil_defaultlib.psb3_0_vector_delay1_x2 
  port map (
    d_1 => slice0_y_net_x0,
    d_2 => slice1_y_net_x0,
    d_3 => slice2_y_net_x0,
    d_4 => slice3_y_net_x0,
    d_5 => slice4_y_net_x0,
    d_6 => slice5_y_net_x0,
    d_7 => slice6_y_net_x0,
    d_8 => slice7_y_net_x0,
    d_9 => slice8_y_net_x0,
    d_10 => slice9_y_net_x0,
    d_11 => slice10_y_net_x0,
    d_12 => slice11_y_net_x0,
    d_13 => slice12_y_net_x0,
    d_14 => slice13_y_net_x0,
    d_15 => slice14_y_net_x0,
    d_16 => slice15_y_net_x0,
    clk_1 => clk_net,
    ce_1 => ce_net,
    q_1 => delay0_q_net,
    q_2 => delay1_q_net,
    q_3 => delay2_q_net,
    q_4 => delay3_q_net,
    q_5 => delay4_q_net,
    q_6 => delay5_q_net,
    q_7 => delay6_q_net,
    q_8 => delay7_q_net,
    q_9 => delay8_q_net,
    q_10 => delay9_q_net,
    q_11 => delay10_q_net,
    q_12 => delay11_q_net,
    q_13 => delay12_q_net,
    q_14 => delay13_q_net,
    q_15 => delay14_q_net,
    q_16 => delay15_q_net
  );
  vector_slice : entity xil_defaultlib.psb3_0_vector_slice_x2 
  port map (
    in_1 => mult0_p_net,
    in_2 => mult1_p_net,
    in_3 => mult2_p_net,
    in_4 => mult3_p_net,
    in_5 => mult4_p_net,
    in_6 => mult5_p_net,
    in_7 => mult6_p_net,
    in_8 => mult7_p_net,
    in_9 => mult8_p_net,
    in_10 => mult9_p_net,
    in_11 => mult10_p_net,
    in_12 => mult11_p_net,
    in_13 => mult12_p_net,
    in_14 => mult13_p_net,
    in_15 => mult14_p_net,
    in_16 => mult15_p_net,
    out_1 => slice0_y_net_x1,
    out_2 => slice1_y_net_x1,
    out_3 => slice2_y_net_x1,
    out_4 => slice3_y_net_x1,
    out_5 => slice4_y_net_x1,
    out_6 => slice5_y_net_x1,
    out_7 => slice6_y_net_x1,
    out_8 => slice7_y_net_x1,
    out_9 => slice8_y_net_x1,
    out_10 => slice9_y_net_x1,
    out_11 => slice10_y_net_x1,
    out_12 => slice11_y_net_x1,
    out_13 => slice12_y_net_x1,
    out_14 => slice13_y_net_x1,
    out_15 => slice14_y_net_x1,
    out_16 => slice15_y_net_x1
  );
  vector_slice1 : entity xil_defaultlib.psb3_0_vector_slice1_x2 
  port map (
    in_1 => reinterpret0_output_port_net,
    in_2 => reinterpret1_output_port_net,
    in_3 => reinterpret2_output_port_net,
    in_4 => reinterpret3_output_port_net,
    in_5 => reinterpret4_output_port_net,
    in_6 => reinterpret5_output_port_net,
    in_7 => reinterpret6_output_port_net,
    in_8 => reinterpret7_output_port_net,
    in_9 => reinterpret8_output_port_net,
    in_10 => reinterpret9_output_port_net,
    in_11 => reinterpret10_output_port_net,
    in_12 => reinterpret11_output_port_net,
    in_13 => reinterpret12_output_port_net,
    in_14 => reinterpret13_output_port_net,
    in_15 => reinterpret14_output_port_net,
    in_16 => reinterpret15_output_port_net,
    out_1 => slice0_y_net_x0,
    out_2 => slice1_y_net_x0,
    out_3 => slice2_y_net_x0,
    out_4 => slice3_y_net_x0,
    out_5 => slice4_y_net_x0,
    out_6 => slice5_y_net_x0,
    out_7 => slice6_y_net_x0,
    out_8 => slice7_y_net_x0,
    out_9 => slice8_y_net_x0,
    out_10 => slice9_y_net_x0,
    out_11 => slice10_y_net_x0,
    out_12 => slice11_y_net_x0,
    out_13 => slice12_y_net_x0,
    out_14 => slice13_y_net_x0,
    out_15 => slice14_y_net_x0,
    out_16 => slice15_y_net_x0
  );
  vector_slice2 : entity xil_defaultlib.psb3_0_vector_slice2_x2 
  port map (
    in_1 => addsub0_s_net,
    in_2 => addsub1_s_net,
    in_3 => addsub2_s_net,
    in_4 => addsub3_s_net,
    in_5 => addsub4_s_net,
    in_6 => addsub5_s_net,
    in_7 => addsub6_s_net,
    in_8 => addsub7_s_net,
    in_9 => addsub8_s_net,
    in_10 => addsub9_s_net,
    in_11 => addsub10_s_net,
    in_12 => addsub11_s_net,
    in_13 => addsub12_s_net,
    in_14 => addsub13_s_net,
    in_15 => addsub14_s_net,
    in_16 => addsub15_s_net,
    out_1 => slice0_y_net,
    out_2 => slice1_y_net,
    out_3 => slice2_y_net,
    out_4 => slice3_y_net,
    out_5 => slice4_y_net,
    out_6 => slice5_y_net,
    out_7 => slice6_y_net,
    out_8 => slice7_y_net,
    out_9 => slice8_y_net,
    out_10 => slice9_y_net,
    out_11 => slice10_y_net,
    out_12 => slice11_y_net,
    out_13 => slice12_y_net,
    out_14 => slice13_y_net,
    out_15 => slice14_y_net,
    out_16 => slice15_y_net
  );
  vector_to_scalar : entity xil_defaultlib.psb3_0_vector_to_scalar_x2 
  port map (
    i_1 => delay0_q_net_x0,
    i_2 => delay1_q_net_x0,
    i_3 => delay2_q_net_x0,
    i_4 => delay3_q_net_x0,
    i_5 => delay4_q_net_x0,
    i_6 => delay5_q_net_x0,
    i_7 => delay6_q_net_x0,
    i_8 => delay7_q_net_x0,
    i_9 => delay8_q_net_x0,
    i_10 => delay9_q_net_x0,
    i_11 => delay10_q_net_x0,
    i_12 => delay11_q_net_x0,
    i_13 => delay12_q_net_x0,
    i_14 => delay13_q_net_x0,
    i_15 => delay14_q_net_x0,
    i_16 => delay15_q_net_x0,
    o => concat1_y_net_x1
  );
  vector_to_scalar1 : entity xil_defaultlib.psb3_0_vector_to_scalar1_x2 
  port map (
    i_1 => delay0_q_net,
    i_2 => delay1_q_net,
    i_3 => delay2_q_net,
    i_4 => delay3_q_net,
    i_5 => delay4_q_net,
    i_6 => delay5_q_net,
    i_7 => delay6_q_net,
    i_8 => delay7_q_net,
    i_9 => delay8_q_net,
    i_10 => delay9_q_net,
    i_11 => delay10_q_net,
    i_12 => delay11_q_net,
    i_13 => delay12_q_net,
    i_14 => delay13_q_net,
    i_15 => delay14_q_net,
    i_16 => delay15_q_net,
    o => concat1_y_net_x0
  );
  vector_to_scalar2 : entity xil_defaultlib.psb3_0_vector_to_scalar2_x2 
  port map (
    i_1 => slice0_y_net,
    i_2 => slice1_y_net,
    i_3 => slice2_y_net,
    i_4 => slice3_y_net,
    i_5 => slice4_y_net,
    i_6 => slice5_y_net,
    i_7 => slice6_y_net,
    i_8 => slice7_y_net,
    i_9 => slice8_y_net,
    i_10 => slice9_y_net,
    i_11 => slice10_y_net,
    i_12 => slice11_y_net,
    i_13 => slice12_y_net,
    i_14 => slice13_y_net,
    i_15 => slice14_y_net,
    i_16 => slice15_y_net,
    o => concat1_y_net
  );
  constant17 : entity xil_defaultlib.sysgen_constant_71e89d757c 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant17_op_net
  );
  convert : entity xil_defaultlib.psb3_0_xlconvert 
  generic map (
    bool_conversion => 1,
    din_arith => 1,
    din_bin_pt => 0,
    din_width => 1,
    dout_arith => 1,
    dout_bin_pt => 0,
    dout_width => 1,
    latency => 1,
    overflow => xlWrap,
    quantization => xlTruncate
  )
  port map (
    clr => '0',
    en => "1",
    din => expression_dout_net,
    clk => clk_net,
    ce => ce_net,
    dout => convert_dout_net
  );
  expression : entity xil_defaultlib.sysgen_expr_7c83532765 
  port map (
    clr => '0',
    a => concat1_y_net_x1,
    b => concat1_y_net_x0,
    s => concat1_y_net,
    clk => clk_net,
    ce => ce_net,
    dout => expression_dout_net
  );
  register_x0 : entity xil_defaultlib.psb3_0_xlregister 
  generic map (
    d_width => 1,
    init_value => b"0"
  )
  port map (
    d => constant17_op_net,
    rst => gin_tl_reset_net,
    en => convert_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => register_q_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Overflow Detector add_re_1/Vector Delay
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_delay_x3 is
  port (
    d_1 : in std_logic_vector( 1-1 downto 0 );
    d_2 : in std_logic_vector( 1-1 downto 0 );
    d_3 : in std_logic_vector( 1-1 downto 0 );
    d_4 : in std_logic_vector( 1-1 downto 0 );
    d_5 : in std_logic_vector( 1-1 downto 0 );
    d_6 : in std_logic_vector( 1-1 downto 0 );
    d_7 : in std_logic_vector( 1-1 downto 0 );
    d_8 : in std_logic_vector( 1-1 downto 0 );
    d_9 : in std_logic_vector( 1-1 downto 0 );
    d_10 : in std_logic_vector( 1-1 downto 0 );
    d_11 : in std_logic_vector( 1-1 downto 0 );
    d_12 : in std_logic_vector( 1-1 downto 0 );
    d_13 : in std_logic_vector( 1-1 downto 0 );
    d_14 : in std_logic_vector( 1-1 downto 0 );
    d_15 : in std_logic_vector( 1-1 downto 0 );
    d_16 : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    q_1 : out std_logic_vector( 1-1 downto 0 );
    q_2 : out std_logic_vector( 1-1 downto 0 );
    q_3 : out std_logic_vector( 1-1 downto 0 );
    q_4 : out std_logic_vector( 1-1 downto 0 );
    q_5 : out std_logic_vector( 1-1 downto 0 );
    q_6 : out std_logic_vector( 1-1 downto 0 );
    q_7 : out std_logic_vector( 1-1 downto 0 );
    q_8 : out std_logic_vector( 1-1 downto 0 );
    q_9 : out std_logic_vector( 1-1 downto 0 );
    q_10 : out std_logic_vector( 1-1 downto 0 );
    q_11 : out std_logic_vector( 1-1 downto 0 );
    q_12 : out std_logic_vector( 1-1 downto 0 );
    q_13 : out std_logic_vector( 1-1 downto 0 );
    q_14 : out std_logic_vector( 1-1 downto 0 );
    q_15 : out std_logic_vector( 1-1 downto 0 );
    q_16 : out std_logic_vector( 1-1 downto 0 )
  );
end psb3_0_vector_delay_x3;
architecture structural of psb3_0_vector_delay_x3 is 
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay12_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay14_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay7_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay0_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay10_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay13_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay9_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay15_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay11_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal slice10_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal slice15_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 1-1 downto 0 );
begin
  q_1 <= delay0_q_net;
  q_2 <= delay1_q_net;
  q_3 <= delay2_q_net;
  q_4 <= delay3_q_net;
  q_5 <= delay4_q_net;
  q_6 <= delay5_q_net;
  q_7 <= delay6_q_net;
  q_8 <= delay7_q_net;
  q_9 <= delay8_q_net;
  q_10 <= delay9_q_net;
  q_11 <= delay10_q_net;
  q_12 <= delay11_q_net;
  q_13 <= delay12_q_net;
  q_14 <= delay13_q_net;
  q_15 <= delay14_q_net;
  q_16 <= delay15_q_net;
  slice0_y_net <= d_1;
  slice1_y_net <= d_2;
  slice2_y_net <= d_3;
  slice3_y_net <= d_4;
  slice4_y_net <= d_5;
  slice5_y_net <= d_6;
  slice6_y_net <= d_7;
  slice7_y_net <= d_8;
  slice8_y_net <= d_9;
  slice9_y_net <= d_10;
  slice10_y_net <= d_11;
  slice11_y_net <= d_12;
  slice12_y_net <= d_13;
  slice13_y_net <= d_14;
  slice14_y_net <= d_15;
  slice15_y_net <= d_16;
  clk_net <= clk_1;
  ce_net <= ce_1;
  delay0 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice0_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay0_q_net
  );
  delay1 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice2_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay3 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice3_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  delay4 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice4_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net
  );
  delay5 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice5_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  delay6 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice6_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay6_q_net
  );
  delay7 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice7_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay7_q_net
  );
  delay8 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice8_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay8_q_net
  );
  delay9 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice9_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay9_q_net
  );
  delay10 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice10_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay10_q_net
  );
  delay11 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice11_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay11_q_net
  );
  delay12 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice12_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay12_q_net
  );
  delay13 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice13_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay13_q_net
  );
  delay14 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice14_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay14_q_net
  );
  delay15 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice15_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay15_q_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Overflow Detector add_re_1/Vector Delay1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_delay1_x3 is
  port (
    d_1 : in std_logic_vector( 1-1 downto 0 );
    d_2 : in std_logic_vector( 1-1 downto 0 );
    d_3 : in std_logic_vector( 1-1 downto 0 );
    d_4 : in std_logic_vector( 1-1 downto 0 );
    d_5 : in std_logic_vector( 1-1 downto 0 );
    d_6 : in std_logic_vector( 1-1 downto 0 );
    d_7 : in std_logic_vector( 1-1 downto 0 );
    d_8 : in std_logic_vector( 1-1 downto 0 );
    d_9 : in std_logic_vector( 1-1 downto 0 );
    d_10 : in std_logic_vector( 1-1 downto 0 );
    d_11 : in std_logic_vector( 1-1 downto 0 );
    d_12 : in std_logic_vector( 1-1 downto 0 );
    d_13 : in std_logic_vector( 1-1 downto 0 );
    d_14 : in std_logic_vector( 1-1 downto 0 );
    d_15 : in std_logic_vector( 1-1 downto 0 );
    d_16 : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    q_1 : out std_logic_vector( 1-1 downto 0 );
    q_2 : out std_logic_vector( 1-1 downto 0 );
    q_3 : out std_logic_vector( 1-1 downto 0 );
    q_4 : out std_logic_vector( 1-1 downto 0 );
    q_5 : out std_logic_vector( 1-1 downto 0 );
    q_6 : out std_logic_vector( 1-1 downto 0 );
    q_7 : out std_logic_vector( 1-1 downto 0 );
    q_8 : out std_logic_vector( 1-1 downto 0 );
    q_9 : out std_logic_vector( 1-1 downto 0 );
    q_10 : out std_logic_vector( 1-1 downto 0 );
    q_11 : out std_logic_vector( 1-1 downto 0 );
    q_12 : out std_logic_vector( 1-1 downto 0 );
    q_13 : out std_logic_vector( 1-1 downto 0 );
    q_14 : out std_logic_vector( 1-1 downto 0 );
    q_15 : out std_logic_vector( 1-1 downto 0 );
    q_16 : out std_logic_vector( 1-1 downto 0 )
  );
end psb3_0_vector_delay1_x3;
architecture structural of psb3_0_vector_delay1_x3 is 
  signal delay0_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay11_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay13_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay9_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay10_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay7_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal slice7_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay12_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay14_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay15_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal slice5_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 1-1 downto 0 );
begin
  q_1 <= delay0_q_net;
  q_2 <= delay1_q_net;
  q_3 <= delay2_q_net;
  q_4 <= delay3_q_net;
  q_5 <= delay4_q_net;
  q_6 <= delay5_q_net;
  q_7 <= delay6_q_net;
  q_8 <= delay7_q_net;
  q_9 <= delay8_q_net;
  q_10 <= delay9_q_net;
  q_11 <= delay10_q_net;
  q_12 <= delay11_q_net;
  q_13 <= delay12_q_net;
  q_14 <= delay13_q_net;
  q_15 <= delay14_q_net;
  q_16 <= delay15_q_net;
  slice0_y_net <= d_1;
  slice1_y_net <= d_2;
  slice2_y_net <= d_3;
  slice3_y_net <= d_4;
  slice4_y_net <= d_5;
  slice5_y_net <= d_6;
  slice6_y_net <= d_7;
  slice7_y_net <= d_8;
  slice8_y_net <= d_9;
  slice9_y_net <= d_10;
  slice10_y_net <= d_11;
  slice11_y_net <= d_12;
  slice12_y_net <= d_13;
  slice13_y_net <= d_14;
  slice14_y_net <= d_15;
  slice15_y_net <= d_16;
  clk_net <= clk_1;
  ce_net <= ce_1;
  delay0 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice0_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay0_q_net
  );
  delay1 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice2_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay3 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice3_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  delay4 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice4_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net
  );
  delay5 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice5_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  delay6 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice6_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay6_q_net
  );
  delay7 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice7_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay7_q_net
  );
  delay8 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice8_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay8_q_net
  );
  delay9 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice9_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay9_q_net
  );
  delay10 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice10_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay10_q_net
  );
  delay11 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice11_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay11_q_net
  );
  delay12 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice12_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay12_q_net
  );
  delay13 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice13_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay13_q_net
  );
  delay14 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice14_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay14_q_net
  );
  delay15 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice15_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay15_q_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Overflow Detector add_re_1/Vector Slice
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_slice_x3 is
  port (
    in_1 : in std_logic_vector( 16-1 downto 0 );
    in_2 : in std_logic_vector( 16-1 downto 0 );
    in_3 : in std_logic_vector( 16-1 downto 0 );
    in_4 : in std_logic_vector( 16-1 downto 0 );
    in_5 : in std_logic_vector( 16-1 downto 0 );
    in_6 : in std_logic_vector( 16-1 downto 0 );
    in_7 : in std_logic_vector( 16-1 downto 0 );
    in_8 : in std_logic_vector( 16-1 downto 0 );
    in_9 : in std_logic_vector( 16-1 downto 0 );
    in_10 : in std_logic_vector( 16-1 downto 0 );
    in_11 : in std_logic_vector( 16-1 downto 0 );
    in_12 : in std_logic_vector( 16-1 downto 0 );
    in_13 : in std_logic_vector( 16-1 downto 0 );
    in_14 : in std_logic_vector( 16-1 downto 0 );
    in_15 : in std_logic_vector( 16-1 downto 0 );
    in_16 : in std_logic_vector( 16-1 downto 0 );
    out_1 : out std_logic_vector( 1-1 downto 0 );
    out_2 : out std_logic_vector( 1-1 downto 0 );
    out_3 : out std_logic_vector( 1-1 downto 0 );
    out_4 : out std_logic_vector( 1-1 downto 0 );
    out_5 : out std_logic_vector( 1-1 downto 0 );
    out_6 : out std_logic_vector( 1-1 downto 0 );
    out_7 : out std_logic_vector( 1-1 downto 0 );
    out_8 : out std_logic_vector( 1-1 downto 0 );
    out_9 : out std_logic_vector( 1-1 downto 0 );
    out_10 : out std_logic_vector( 1-1 downto 0 );
    out_11 : out std_logic_vector( 1-1 downto 0 );
    out_12 : out std_logic_vector( 1-1 downto 0 );
    out_13 : out std_logic_vector( 1-1 downto 0 );
    out_14 : out std_logic_vector( 1-1 downto 0 );
    out_15 : out std_logic_vector( 1-1 downto 0 );
    out_16 : out std_logic_vector( 1-1 downto 0 )
  );
end psb3_0_vector_slice_x3;
architecture structural of psb3_0_vector_slice_x3 is 
  signal slice1_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 1-1 downto 0 );
  signal mult0_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult1_p_net : std_logic_vector( 16-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 1-1 downto 0 );
  signal mult2_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult3_p_net : std_logic_vector( 16-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 1-1 downto 0 );
  signal mult11_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult9_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult13_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult6_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult15_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult8_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult4_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult7_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult12_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult10_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult5_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult14_p_net : std_logic_vector( 16-1 downto 0 );
begin
  out_1 <= slice0_y_net;
  out_2 <= slice1_y_net;
  out_3 <= slice2_y_net;
  out_4 <= slice3_y_net;
  out_5 <= slice4_y_net;
  out_6 <= slice5_y_net;
  out_7 <= slice6_y_net;
  out_8 <= slice7_y_net;
  out_9 <= slice8_y_net;
  out_10 <= slice9_y_net;
  out_11 <= slice10_y_net;
  out_12 <= slice11_y_net;
  out_13 <= slice12_y_net;
  out_14 <= slice13_y_net;
  out_15 <= slice14_y_net;
  out_16 <= slice15_y_net;
  mult0_p_net <= in_1;
  mult1_p_net <= in_2;
  mult2_p_net <= in_3;
  mult3_p_net <= in_4;
  mult4_p_net <= in_5;
  mult5_p_net <= in_6;
  mult6_p_net <= in_7;
  mult7_p_net <= in_8;
  mult8_p_net <= in_9;
  mult9_p_net <= in_10;
  mult10_p_net <= in_11;
  mult11_p_net <= in_12;
  mult12_p_net <= in_13;
  mult13_p_net <= in_14;
  mult14_p_net <= in_15;
  mult15_p_net <= in_16;
  slice0 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult0_p_net,
    y => slice0_y_net
  );
  slice1 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult1_p_net,
    y => slice1_y_net
  );
  slice2 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult2_p_net,
    y => slice2_y_net
  );
  slice3 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult3_p_net,
    y => slice3_y_net
  );
  slice4 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult4_p_net,
    y => slice4_y_net
  );
  slice5 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult5_p_net,
    y => slice5_y_net
  );
  slice6 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult6_p_net,
    y => slice6_y_net
  );
  slice7 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult7_p_net,
    y => slice7_y_net
  );
  slice8 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult8_p_net,
    y => slice8_y_net
  );
  slice9 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult9_p_net,
    y => slice9_y_net
  );
  slice10 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult10_p_net,
    y => slice10_y_net
  );
  slice11 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult11_p_net,
    y => slice11_y_net
  );
  slice12 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult12_p_net,
    y => slice12_y_net
  );
  slice13 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult13_p_net,
    y => slice13_y_net
  );
  slice14 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult14_p_net,
    y => slice14_y_net
  );
  slice15 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult15_p_net,
    y => slice15_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Overflow Detector add_re_1/Vector Slice1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_slice1_x3 is
  port (
    in_1 : in std_logic_vector( 16-1 downto 0 );
    in_2 : in std_logic_vector( 16-1 downto 0 );
    in_3 : in std_logic_vector( 16-1 downto 0 );
    in_4 : in std_logic_vector( 16-1 downto 0 );
    in_5 : in std_logic_vector( 16-1 downto 0 );
    in_6 : in std_logic_vector( 16-1 downto 0 );
    in_7 : in std_logic_vector( 16-1 downto 0 );
    in_8 : in std_logic_vector( 16-1 downto 0 );
    in_9 : in std_logic_vector( 16-1 downto 0 );
    in_10 : in std_logic_vector( 16-1 downto 0 );
    in_11 : in std_logic_vector( 16-1 downto 0 );
    in_12 : in std_logic_vector( 16-1 downto 0 );
    in_13 : in std_logic_vector( 16-1 downto 0 );
    in_14 : in std_logic_vector( 16-1 downto 0 );
    in_15 : in std_logic_vector( 16-1 downto 0 );
    in_16 : in std_logic_vector( 16-1 downto 0 );
    out_1 : out std_logic_vector( 1-1 downto 0 );
    out_2 : out std_logic_vector( 1-1 downto 0 );
    out_3 : out std_logic_vector( 1-1 downto 0 );
    out_4 : out std_logic_vector( 1-1 downto 0 );
    out_5 : out std_logic_vector( 1-1 downto 0 );
    out_6 : out std_logic_vector( 1-1 downto 0 );
    out_7 : out std_logic_vector( 1-1 downto 0 );
    out_8 : out std_logic_vector( 1-1 downto 0 );
    out_9 : out std_logic_vector( 1-1 downto 0 );
    out_10 : out std_logic_vector( 1-1 downto 0 );
    out_11 : out std_logic_vector( 1-1 downto 0 );
    out_12 : out std_logic_vector( 1-1 downto 0 );
    out_13 : out std_logic_vector( 1-1 downto 0 );
    out_14 : out std_logic_vector( 1-1 downto 0 );
    out_15 : out std_logic_vector( 1-1 downto 0 );
    out_16 : out std_logic_vector( 1-1 downto 0 )
  );
end psb3_0_vector_slice1_x3;
architecture structural of psb3_0_vector_slice1_x3 is 
  signal slice3_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
begin
  out_1 <= slice0_y_net;
  out_2 <= slice1_y_net;
  out_3 <= slice2_y_net;
  out_4 <= slice3_y_net;
  out_5 <= slice4_y_net;
  out_6 <= slice5_y_net;
  out_7 <= slice6_y_net;
  out_8 <= slice7_y_net;
  out_9 <= slice8_y_net;
  out_10 <= slice9_y_net;
  out_11 <= slice10_y_net;
  out_12 <= slice11_y_net;
  out_13 <= slice12_y_net;
  out_14 <= slice13_y_net;
  out_15 <= slice14_y_net;
  out_16 <= slice15_y_net;
  reinterpret0_output_port_net <= in_1;
  reinterpret1_output_port_net <= in_2;
  reinterpret2_output_port_net <= in_3;
  reinterpret3_output_port_net <= in_4;
  reinterpret4_output_port_net <= in_5;
  reinterpret5_output_port_net <= in_6;
  reinterpret6_output_port_net <= in_7;
  reinterpret7_output_port_net <= in_8;
  reinterpret8_output_port_net <= in_9;
  reinterpret9_output_port_net <= in_10;
  reinterpret10_output_port_net <= in_11;
  reinterpret11_output_port_net <= in_12;
  reinterpret12_output_port_net <= in_13;
  reinterpret13_output_port_net <= in_14;
  reinterpret14_output_port_net <= in_15;
  reinterpret15_output_port_net <= in_16;
  slice0 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret0_output_port_net,
    y => slice0_y_net
  );
  slice1 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret1_output_port_net,
    y => slice1_y_net
  );
  slice2 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret2_output_port_net,
    y => slice2_y_net
  );
  slice3 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret3_output_port_net,
    y => slice3_y_net
  );
  slice4 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret4_output_port_net,
    y => slice4_y_net
  );
  slice5 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret5_output_port_net,
    y => slice5_y_net
  );
  slice6 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret6_output_port_net,
    y => slice6_y_net
  );
  slice7 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret7_output_port_net,
    y => slice7_y_net
  );
  slice8 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret8_output_port_net,
    y => slice8_y_net
  );
  slice9 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret9_output_port_net,
    y => slice9_y_net
  );
  slice10 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret10_output_port_net,
    y => slice10_y_net
  );
  slice11 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret11_output_port_net,
    y => slice11_y_net
  );
  slice12 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret12_output_port_net,
    y => slice12_y_net
  );
  slice13 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret13_output_port_net,
    y => slice13_y_net
  );
  slice14 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret14_output_port_net,
    y => slice14_y_net
  );
  slice15 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret15_output_port_net,
    y => slice15_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Overflow Detector add_re_1/Vector Slice2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_slice2_x3 is
  port (
    in_1 : in std_logic_vector( 16-1 downto 0 );
    in_2 : in std_logic_vector( 16-1 downto 0 );
    in_3 : in std_logic_vector( 16-1 downto 0 );
    in_4 : in std_logic_vector( 16-1 downto 0 );
    in_5 : in std_logic_vector( 16-1 downto 0 );
    in_6 : in std_logic_vector( 16-1 downto 0 );
    in_7 : in std_logic_vector( 16-1 downto 0 );
    in_8 : in std_logic_vector( 16-1 downto 0 );
    in_9 : in std_logic_vector( 16-1 downto 0 );
    in_10 : in std_logic_vector( 16-1 downto 0 );
    in_11 : in std_logic_vector( 16-1 downto 0 );
    in_12 : in std_logic_vector( 16-1 downto 0 );
    in_13 : in std_logic_vector( 16-1 downto 0 );
    in_14 : in std_logic_vector( 16-1 downto 0 );
    in_15 : in std_logic_vector( 16-1 downto 0 );
    in_16 : in std_logic_vector( 16-1 downto 0 );
    out_1 : out std_logic_vector( 1-1 downto 0 );
    out_2 : out std_logic_vector( 1-1 downto 0 );
    out_3 : out std_logic_vector( 1-1 downto 0 );
    out_4 : out std_logic_vector( 1-1 downto 0 );
    out_5 : out std_logic_vector( 1-1 downto 0 );
    out_6 : out std_logic_vector( 1-1 downto 0 );
    out_7 : out std_logic_vector( 1-1 downto 0 );
    out_8 : out std_logic_vector( 1-1 downto 0 );
    out_9 : out std_logic_vector( 1-1 downto 0 );
    out_10 : out std_logic_vector( 1-1 downto 0 );
    out_11 : out std_logic_vector( 1-1 downto 0 );
    out_12 : out std_logic_vector( 1-1 downto 0 );
    out_13 : out std_logic_vector( 1-1 downto 0 );
    out_14 : out std_logic_vector( 1-1 downto 0 );
    out_15 : out std_logic_vector( 1-1 downto 0 );
    out_16 : out std_logic_vector( 1-1 downto 0 )
  );
end psb3_0_vector_slice2_x3;
architecture structural of psb3_0_vector_slice2_x3 is 
  signal addsub0_s_net : std_logic_vector( 16-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 1-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 16-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 1-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 16-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 1-1 downto 0 );
  signal addsub14_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub15_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub13_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub10_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub3_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub11_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub7_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub9_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub12_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub6_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub5_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub8_s_net : std_logic_vector( 16-1 downto 0 );
begin
  out_1 <= slice0_y_net;
  out_2 <= slice1_y_net;
  out_3 <= slice2_y_net;
  out_4 <= slice3_y_net;
  out_5 <= slice4_y_net;
  out_6 <= slice5_y_net;
  out_7 <= slice6_y_net;
  out_8 <= slice7_y_net;
  out_9 <= slice8_y_net;
  out_10 <= slice9_y_net;
  out_11 <= slice10_y_net;
  out_12 <= slice11_y_net;
  out_13 <= slice12_y_net;
  out_14 <= slice13_y_net;
  out_15 <= slice14_y_net;
  out_16 <= slice15_y_net;
  addsub0_s_net <= in_1;
  addsub1_s_net <= in_2;
  addsub2_s_net <= in_3;
  addsub3_s_net <= in_4;
  addsub4_s_net <= in_5;
  addsub5_s_net <= in_6;
  addsub6_s_net <= in_7;
  addsub7_s_net <= in_8;
  addsub8_s_net <= in_9;
  addsub9_s_net <= in_10;
  addsub10_s_net <= in_11;
  addsub11_s_net <= in_12;
  addsub12_s_net <= in_13;
  addsub13_s_net <= in_14;
  addsub14_s_net <= in_15;
  addsub15_s_net <= in_16;
  slice0 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub0_s_net,
    y => slice0_y_net
  );
  slice1 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub1_s_net,
    y => slice1_y_net
  );
  slice2 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub2_s_net,
    y => slice2_y_net
  );
  slice3 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub3_s_net,
    y => slice3_y_net
  );
  slice4 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub4_s_net,
    y => slice4_y_net
  );
  slice5 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub5_s_net,
    y => slice5_y_net
  );
  slice6 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub6_s_net,
    y => slice6_y_net
  );
  slice7 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub7_s_net,
    y => slice7_y_net
  );
  slice8 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub8_s_net,
    y => slice8_y_net
  );
  slice9 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub9_s_net,
    y => slice9_y_net
  );
  slice10 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub10_s_net,
    y => slice10_y_net
  );
  slice11 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub11_s_net,
    y => slice11_y_net
  );
  slice12 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub12_s_net,
    y => slice12_y_net
  );
  slice13 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub13_s_net,
    y => slice13_y_net
  );
  slice14 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub14_s_net,
    y => slice14_y_net
  );
  slice15 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub15_s_net,
    y => slice15_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Overflow Detector add_re_1/Vector to Scalar
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_to_scalar_x3 is
  port (
    i_1 : in std_logic_vector( 1-1 downto 0 );
    i_2 : in std_logic_vector( 1-1 downto 0 );
    i_3 : in std_logic_vector( 1-1 downto 0 );
    i_4 : in std_logic_vector( 1-1 downto 0 );
    i_5 : in std_logic_vector( 1-1 downto 0 );
    i_6 : in std_logic_vector( 1-1 downto 0 );
    i_7 : in std_logic_vector( 1-1 downto 0 );
    i_8 : in std_logic_vector( 1-1 downto 0 );
    i_9 : in std_logic_vector( 1-1 downto 0 );
    i_10 : in std_logic_vector( 1-1 downto 0 );
    i_11 : in std_logic_vector( 1-1 downto 0 );
    i_12 : in std_logic_vector( 1-1 downto 0 );
    i_13 : in std_logic_vector( 1-1 downto 0 );
    i_14 : in std_logic_vector( 1-1 downto 0 );
    i_15 : in std_logic_vector( 1-1 downto 0 );
    i_16 : in std_logic_vector( 1-1 downto 0 );
    o : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_vector_to_scalar_x3;
architecture structural of psb3_0_vector_to_scalar_x3 is 
  signal concat1_y_net : std_logic_vector( 16-1 downto 0 );
  signal delay0_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay13_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay11_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay7_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay9_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay15_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay12_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay10_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay14_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 1-1 downto 0 );
begin
  o <= concat1_y_net;
  delay0_q_net <= i_1;
  delay1_q_net <= i_2;
  delay2_q_net <= i_3;
  delay3_q_net <= i_4;
  delay4_q_net <= i_5;
  delay5_q_net <= i_6;
  delay6_q_net <= i_7;
  delay7_q_net <= i_8;
  delay8_q_net <= i_9;
  delay9_q_net <= i_10;
  delay10_q_net <= i_11;
  delay11_q_net <= i_12;
  delay12_q_net <= i_13;
  delay13_q_net <= i_14;
  delay14_q_net <= i_15;
  delay15_q_net <= i_16;
  concat1 : entity xil_defaultlib.sysgen_concat_d977c66e35 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => delay15_q_net,
    in1 => delay14_q_net,
    in2 => delay13_q_net,
    in3 => delay12_q_net,
    in4 => delay11_q_net,
    in5 => delay10_q_net,
    in6 => delay9_q_net,
    in7 => delay8_q_net,
    in8 => delay7_q_net,
    in9 => delay6_q_net,
    in10 => delay5_q_net,
    in11 => delay4_q_net,
    in12 => delay3_q_net,
    in13 => delay2_q_net,
    in14 => delay1_q_net,
    in15 => delay0_q_net,
    y => concat1_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Overflow Detector add_re_1/Vector to Scalar1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_to_scalar1_x3 is
  port (
    i_1 : in std_logic_vector( 1-1 downto 0 );
    i_2 : in std_logic_vector( 1-1 downto 0 );
    i_3 : in std_logic_vector( 1-1 downto 0 );
    i_4 : in std_logic_vector( 1-1 downto 0 );
    i_5 : in std_logic_vector( 1-1 downto 0 );
    i_6 : in std_logic_vector( 1-1 downto 0 );
    i_7 : in std_logic_vector( 1-1 downto 0 );
    i_8 : in std_logic_vector( 1-1 downto 0 );
    i_9 : in std_logic_vector( 1-1 downto 0 );
    i_10 : in std_logic_vector( 1-1 downto 0 );
    i_11 : in std_logic_vector( 1-1 downto 0 );
    i_12 : in std_logic_vector( 1-1 downto 0 );
    i_13 : in std_logic_vector( 1-1 downto 0 );
    i_14 : in std_logic_vector( 1-1 downto 0 );
    i_15 : in std_logic_vector( 1-1 downto 0 );
    i_16 : in std_logic_vector( 1-1 downto 0 );
    o : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_vector_to_scalar1_x3;
architecture structural of psb3_0_vector_to_scalar1_x3 is 
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 1-1 downto 0 );
  signal concat1_y_net : std_logic_vector( 16-1 downto 0 );
  signal delay0_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay11_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay12_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay14_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay13_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay9_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay7_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay10_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay15_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
begin
  o <= concat1_y_net;
  delay0_q_net <= i_1;
  delay1_q_net <= i_2;
  delay2_q_net <= i_3;
  delay3_q_net <= i_4;
  delay4_q_net <= i_5;
  delay5_q_net <= i_6;
  delay6_q_net <= i_7;
  delay7_q_net <= i_8;
  delay8_q_net <= i_9;
  delay9_q_net <= i_10;
  delay10_q_net <= i_11;
  delay11_q_net <= i_12;
  delay12_q_net <= i_13;
  delay13_q_net <= i_14;
  delay14_q_net <= i_15;
  delay15_q_net <= i_16;
  concat1 : entity xil_defaultlib.sysgen_concat_d977c66e35 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => delay15_q_net,
    in1 => delay14_q_net,
    in2 => delay13_q_net,
    in3 => delay12_q_net,
    in4 => delay11_q_net,
    in5 => delay10_q_net,
    in6 => delay9_q_net,
    in7 => delay8_q_net,
    in8 => delay7_q_net,
    in9 => delay6_q_net,
    in10 => delay5_q_net,
    in11 => delay4_q_net,
    in12 => delay3_q_net,
    in13 => delay2_q_net,
    in14 => delay1_q_net,
    in15 => delay0_q_net,
    y => concat1_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Overflow Detector add_re_1/Vector to Scalar2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_to_scalar2_x3 is
  port (
    i_1 : in std_logic_vector( 1-1 downto 0 );
    i_2 : in std_logic_vector( 1-1 downto 0 );
    i_3 : in std_logic_vector( 1-1 downto 0 );
    i_4 : in std_logic_vector( 1-1 downto 0 );
    i_5 : in std_logic_vector( 1-1 downto 0 );
    i_6 : in std_logic_vector( 1-1 downto 0 );
    i_7 : in std_logic_vector( 1-1 downto 0 );
    i_8 : in std_logic_vector( 1-1 downto 0 );
    i_9 : in std_logic_vector( 1-1 downto 0 );
    i_10 : in std_logic_vector( 1-1 downto 0 );
    i_11 : in std_logic_vector( 1-1 downto 0 );
    i_12 : in std_logic_vector( 1-1 downto 0 );
    i_13 : in std_logic_vector( 1-1 downto 0 );
    i_14 : in std_logic_vector( 1-1 downto 0 );
    i_15 : in std_logic_vector( 1-1 downto 0 );
    i_16 : in std_logic_vector( 1-1 downto 0 );
    o : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_vector_to_scalar2_x3;
architecture structural of psb3_0_vector_to_scalar2_x3 is 
  signal slice3_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 1-1 downto 0 );
  signal concat1_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 1-1 downto 0 );
begin
  o <= concat1_y_net;
  slice0_y_net <= i_1;
  slice1_y_net <= i_2;
  slice2_y_net <= i_3;
  slice3_y_net <= i_4;
  slice4_y_net <= i_5;
  slice5_y_net <= i_6;
  slice6_y_net <= i_7;
  slice7_y_net <= i_8;
  slice8_y_net <= i_9;
  slice9_y_net <= i_10;
  slice10_y_net <= i_11;
  slice11_y_net <= i_12;
  slice12_y_net <= i_13;
  slice13_y_net <= i_14;
  slice14_y_net <= i_15;
  slice15_y_net <= i_16;
  concat1 : entity xil_defaultlib.sysgen_concat_d977c66e35 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => slice15_y_net,
    in1 => slice14_y_net,
    in2 => slice13_y_net,
    in3 => slice12_y_net,
    in4 => slice11_y_net,
    in5 => slice10_y_net,
    in6 => slice9_y_net,
    in7 => slice8_y_net,
    in8 => slice7_y_net,
    in9 => slice6_y_net,
    in10 => slice5_y_net,
    in11 => slice4_y_net,
    in12 => slice3_y_net,
    in13 => slice2_y_net,
    in14 => slice1_y_net,
    in15 => slice0_y_net,
    y => concat1_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Overflow Detector add_re_1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_overflow_detector_add_re_1 is
  port (
    rst : in std_logic_vector( 1-1 downto 0 );
    a_1 : in std_logic_vector( 16-1 downto 0 );
    b_1 : in std_logic_vector( 16-1 downto 0 );
    s_1 : in std_logic_vector( 16-1 downto 0 );
    a_2 : in std_logic_vector( 16-1 downto 0 );
    a_3 : in std_logic_vector( 16-1 downto 0 );
    a_4 : in std_logic_vector( 16-1 downto 0 );
    a_5 : in std_logic_vector( 16-1 downto 0 );
    a_6 : in std_logic_vector( 16-1 downto 0 );
    a_7 : in std_logic_vector( 16-1 downto 0 );
    a_8 : in std_logic_vector( 16-1 downto 0 );
    a_9 : in std_logic_vector( 16-1 downto 0 );
    a_10 : in std_logic_vector( 16-1 downto 0 );
    a_11 : in std_logic_vector( 16-1 downto 0 );
    a_12 : in std_logic_vector( 16-1 downto 0 );
    a_13 : in std_logic_vector( 16-1 downto 0 );
    a_14 : in std_logic_vector( 16-1 downto 0 );
    a_15 : in std_logic_vector( 16-1 downto 0 );
    a_16 : in std_logic_vector( 16-1 downto 0 );
    b_2 : in std_logic_vector( 16-1 downto 0 );
    b_3 : in std_logic_vector( 16-1 downto 0 );
    b_4 : in std_logic_vector( 16-1 downto 0 );
    b_5 : in std_logic_vector( 16-1 downto 0 );
    b_6 : in std_logic_vector( 16-1 downto 0 );
    b_7 : in std_logic_vector( 16-1 downto 0 );
    b_8 : in std_logic_vector( 16-1 downto 0 );
    b_9 : in std_logic_vector( 16-1 downto 0 );
    b_10 : in std_logic_vector( 16-1 downto 0 );
    b_11 : in std_logic_vector( 16-1 downto 0 );
    b_12 : in std_logic_vector( 16-1 downto 0 );
    b_13 : in std_logic_vector( 16-1 downto 0 );
    b_14 : in std_logic_vector( 16-1 downto 0 );
    b_15 : in std_logic_vector( 16-1 downto 0 );
    b_16 : in std_logic_vector( 16-1 downto 0 );
    s_2 : in std_logic_vector( 16-1 downto 0 );
    s_3 : in std_logic_vector( 16-1 downto 0 );
    s_4 : in std_logic_vector( 16-1 downto 0 );
    s_5 : in std_logic_vector( 16-1 downto 0 );
    s_6 : in std_logic_vector( 16-1 downto 0 );
    s_7 : in std_logic_vector( 16-1 downto 0 );
    s_8 : in std_logic_vector( 16-1 downto 0 );
    s_9 : in std_logic_vector( 16-1 downto 0 );
    s_10 : in std_logic_vector( 16-1 downto 0 );
    s_11 : in std_logic_vector( 16-1 downto 0 );
    s_12 : in std_logic_vector( 16-1 downto 0 );
    s_13 : in std_logic_vector( 16-1 downto 0 );
    s_14 : in std_logic_vector( 16-1 downto 0 );
    s_15 : in std_logic_vector( 16-1 downto 0 );
    s_16 : in std_logic_vector( 16-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    ov : out std_logic_vector( 1-1 downto 0 )
  );
end psb3_0_overflow_detector_add_re_1;
architecture structural of psb3_0_overflow_detector_add_re_1 is 
  signal mult6_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult7_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult9_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult0_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult8_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult3_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult10_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult11_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult4_p_net : std_logic_vector( 16-1 downto 0 );
  signal addsub0_s_net : std_logic_vector( 16-1 downto 0 );
  signal register_q_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mult1_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult2_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult5_p_net : std_logic_vector( 16-1 downto 0 );
  signal gin_tl_reset_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mult12_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult13_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub5_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub3_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub7_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub10_s_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub13_s_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mult14_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mult15_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub6_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub8_s_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub9_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub11_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub12_s_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 16-1 downto 0 );
  signal delay13_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice1_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay4_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay15_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice11_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay15_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice3_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice4_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice5_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice6_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay12_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice13_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal slice7_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice8_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal delay10_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal delay3_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice8_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay5_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay0_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice3_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice7_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 1-1 downto 0 );
  signal addsub14_s_net : std_logic_vector( 16-1 downto 0 );
  signal delay14_q_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal addsub15_s_net : std_logic_vector( 16-1 downto 0 );
  signal delay6_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay7_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice0_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal slice2_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal delay12_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice15_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay14_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay13_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice6_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal delay10_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay8_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay9_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay11_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice5_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal delay7_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice0_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice1_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal slice12_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice2_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice4_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal slice10_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal slice14_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal delay0_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay11_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice9_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal delay9_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice14_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice9_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 1-1 downto 0 );
  signal concat1_y_net_x1 : std_logic_vector( 16-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice13_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 1-1 downto 0 );
  signal constant17_op_net : std_logic_vector( 1-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 1-1 downto 0 );
  signal concat1_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 1-1 downto 0 );
  signal expression_dout_net : std_logic_vector( 1-1 downto 0 );
  signal slice10_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 1-1 downto 0 );
  signal concat1_y_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice15_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal convert_dout_net : std_logic_vector( 1-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice12_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice11_y_net_x0 : std_logic_vector( 1-1 downto 0 );
begin
  ov <= register_q_net;
  gin_tl_reset_net <= rst;
  mult0_p_net <= a_1;
  reinterpret0_output_port_net <= b_1;
  addsub0_s_net <= s_1;
  mult1_p_net <= a_2;
  mult2_p_net <= a_3;
  mult3_p_net <= a_4;
  mult4_p_net <= a_5;
  mult5_p_net <= a_6;
  mult6_p_net <= a_7;
  mult7_p_net <= a_8;
  mult8_p_net <= a_9;
  mult9_p_net <= a_10;
  mult10_p_net <= a_11;
  mult11_p_net <= a_12;
  mult12_p_net <= a_13;
  mult13_p_net <= a_14;
  mult14_p_net <= a_15;
  mult15_p_net <= a_16;
  reinterpret1_output_port_net <= b_2;
  reinterpret2_output_port_net <= b_3;
  reinterpret3_output_port_net <= b_4;
  reinterpret4_output_port_net <= b_5;
  reinterpret5_output_port_net <= b_6;
  reinterpret6_output_port_net <= b_7;
  reinterpret7_output_port_net <= b_8;
  reinterpret8_output_port_net <= b_9;
  reinterpret9_output_port_net <= b_10;
  reinterpret10_output_port_net <= b_11;
  reinterpret11_output_port_net <= b_12;
  reinterpret12_output_port_net <= b_13;
  reinterpret13_output_port_net <= b_14;
  reinterpret14_output_port_net <= b_15;
  reinterpret15_output_port_net <= b_16;
  addsub1_s_net <= s_2;
  addsub2_s_net <= s_3;
  addsub3_s_net <= s_4;
  addsub4_s_net <= s_5;
  addsub5_s_net <= s_6;
  addsub6_s_net <= s_7;
  addsub7_s_net <= s_8;
  addsub8_s_net <= s_9;
  addsub9_s_net <= s_10;
  addsub10_s_net <= s_11;
  addsub11_s_net <= s_12;
  addsub12_s_net <= s_13;
  addsub13_s_net <= s_14;
  addsub14_s_net <= s_15;
  addsub15_s_net <= s_16;
  clk_net <= clk_1;
  ce_net <= ce_1;
  vector_delay : entity xil_defaultlib.psb3_0_vector_delay_x3 
  port map (
    d_1 => slice0_y_net_x1,
    d_2 => slice1_y_net_x1,
    d_3 => slice2_y_net_x1,
    d_4 => slice3_y_net_x1,
    d_5 => slice4_y_net_x1,
    d_6 => slice5_y_net_x1,
    d_7 => slice6_y_net_x1,
    d_8 => slice7_y_net_x1,
    d_9 => slice8_y_net_x1,
    d_10 => slice9_y_net_x1,
    d_11 => slice10_y_net_x1,
    d_12 => slice11_y_net_x1,
    d_13 => slice12_y_net_x1,
    d_14 => slice13_y_net_x1,
    d_15 => slice14_y_net_x1,
    d_16 => slice15_y_net_x1,
    clk_1 => clk_net,
    ce_1 => ce_net,
    q_1 => delay0_q_net_x0,
    q_2 => delay1_q_net_x0,
    q_3 => delay2_q_net_x0,
    q_4 => delay3_q_net_x0,
    q_5 => delay4_q_net_x0,
    q_6 => delay5_q_net_x0,
    q_7 => delay6_q_net_x0,
    q_8 => delay7_q_net_x0,
    q_9 => delay8_q_net_x0,
    q_10 => delay9_q_net_x0,
    q_11 => delay10_q_net_x0,
    q_12 => delay11_q_net_x0,
    q_13 => delay12_q_net_x0,
    q_14 => delay13_q_net_x0,
    q_15 => delay14_q_net_x0,
    q_16 => delay15_q_net_x0
  );
  vector_delay1 : entity xil_defaultlib.psb3_0_vector_delay1_x3 
  port map (
    d_1 => slice0_y_net_x0,
    d_2 => slice1_y_net_x0,
    d_3 => slice2_y_net_x0,
    d_4 => slice3_y_net_x0,
    d_5 => slice4_y_net_x0,
    d_6 => slice5_y_net_x0,
    d_7 => slice6_y_net_x0,
    d_8 => slice7_y_net_x0,
    d_9 => slice8_y_net_x0,
    d_10 => slice9_y_net_x0,
    d_11 => slice10_y_net_x0,
    d_12 => slice11_y_net_x0,
    d_13 => slice12_y_net_x0,
    d_14 => slice13_y_net_x0,
    d_15 => slice14_y_net_x0,
    d_16 => slice15_y_net_x0,
    clk_1 => clk_net,
    ce_1 => ce_net,
    q_1 => delay0_q_net,
    q_2 => delay1_q_net,
    q_3 => delay2_q_net,
    q_4 => delay3_q_net,
    q_5 => delay4_q_net,
    q_6 => delay5_q_net,
    q_7 => delay6_q_net,
    q_8 => delay7_q_net,
    q_9 => delay8_q_net,
    q_10 => delay9_q_net,
    q_11 => delay10_q_net,
    q_12 => delay11_q_net,
    q_13 => delay12_q_net,
    q_14 => delay13_q_net,
    q_15 => delay14_q_net,
    q_16 => delay15_q_net
  );
  vector_slice : entity xil_defaultlib.psb3_0_vector_slice_x3 
  port map (
    in_1 => mult0_p_net,
    in_2 => mult1_p_net,
    in_3 => mult2_p_net,
    in_4 => mult3_p_net,
    in_5 => mult4_p_net,
    in_6 => mult5_p_net,
    in_7 => mult6_p_net,
    in_8 => mult7_p_net,
    in_9 => mult8_p_net,
    in_10 => mult9_p_net,
    in_11 => mult10_p_net,
    in_12 => mult11_p_net,
    in_13 => mult12_p_net,
    in_14 => mult13_p_net,
    in_15 => mult14_p_net,
    in_16 => mult15_p_net,
    out_1 => slice0_y_net_x1,
    out_2 => slice1_y_net_x1,
    out_3 => slice2_y_net_x1,
    out_4 => slice3_y_net_x1,
    out_5 => slice4_y_net_x1,
    out_6 => slice5_y_net_x1,
    out_7 => slice6_y_net_x1,
    out_8 => slice7_y_net_x1,
    out_9 => slice8_y_net_x1,
    out_10 => slice9_y_net_x1,
    out_11 => slice10_y_net_x1,
    out_12 => slice11_y_net_x1,
    out_13 => slice12_y_net_x1,
    out_14 => slice13_y_net_x1,
    out_15 => slice14_y_net_x1,
    out_16 => slice15_y_net_x1
  );
  vector_slice1 : entity xil_defaultlib.psb3_0_vector_slice1_x3 
  port map (
    in_1 => reinterpret0_output_port_net,
    in_2 => reinterpret1_output_port_net,
    in_3 => reinterpret2_output_port_net,
    in_4 => reinterpret3_output_port_net,
    in_5 => reinterpret4_output_port_net,
    in_6 => reinterpret5_output_port_net,
    in_7 => reinterpret6_output_port_net,
    in_8 => reinterpret7_output_port_net,
    in_9 => reinterpret8_output_port_net,
    in_10 => reinterpret9_output_port_net,
    in_11 => reinterpret10_output_port_net,
    in_12 => reinterpret11_output_port_net,
    in_13 => reinterpret12_output_port_net,
    in_14 => reinterpret13_output_port_net,
    in_15 => reinterpret14_output_port_net,
    in_16 => reinterpret15_output_port_net,
    out_1 => slice0_y_net_x0,
    out_2 => slice1_y_net_x0,
    out_3 => slice2_y_net_x0,
    out_4 => slice3_y_net_x0,
    out_5 => slice4_y_net_x0,
    out_6 => slice5_y_net_x0,
    out_7 => slice6_y_net_x0,
    out_8 => slice7_y_net_x0,
    out_9 => slice8_y_net_x0,
    out_10 => slice9_y_net_x0,
    out_11 => slice10_y_net_x0,
    out_12 => slice11_y_net_x0,
    out_13 => slice12_y_net_x0,
    out_14 => slice13_y_net_x0,
    out_15 => slice14_y_net_x0,
    out_16 => slice15_y_net_x0
  );
  vector_slice2 : entity xil_defaultlib.psb3_0_vector_slice2_x3 
  port map (
    in_1 => addsub0_s_net,
    in_2 => addsub1_s_net,
    in_3 => addsub2_s_net,
    in_4 => addsub3_s_net,
    in_5 => addsub4_s_net,
    in_6 => addsub5_s_net,
    in_7 => addsub6_s_net,
    in_8 => addsub7_s_net,
    in_9 => addsub8_s_net,
    in_10 => addsub9_s_net,
    in_11 => addsub10_s_net,
    in_12 => addsub11_s_net,
    in_13 => addsub12_s_net,
    in_14 => addsub13_s_net,
    in_15 => addsub14_s_net,
    in_16 => addsub15_s_net,
    out_1 => slice0_y_net,
    out_2 => slice1_y_net,
    out_3 => slice2_y_net,
    out_4 => slice3_y_net,
    out_5 => slice4_y_net,
    out_6 => slice5_y_net,
    out_7 => slice6_y_net,
    out_8 => slice7_y_net,
    out_9 => slice8_y_net,
    out_10 => slice9_y_net,
    out_11 => slice10_y_net,
    out_12 => slice11_y_net,
    out_13 => slice12_y_net,
    out_14 => slice13_y_net,
    out_15 => slice14_y_net,
    out_16 => slice15_y_net
  );
  vector_to_scalar : entity xil_defaultlib.psb3_0_vector_to_scalar_x3 
  port map (
    i_1 => delay0_q_net_x0,
    i_2 => delay1_q_net_x0,
    i_3 => delay2_q_net_x0,
    i_4 => delay3_q_net_x0,
    i_5 => delay4_q_net_x0,
    i_6 => delay5_q_net_x0,
    i_7 => delay6_q_net_x0,
    i_8 => delay7_q_net_x0,
    i_9 => delay8_q_net_x0,
    i_10 => delay9_q_net_x0,
    i_11 => delay10_q_net_x0,
    i_12 => delay11_q_net_x0,
    i_13 => delay12_q_net_x0,
    i_14 => delay13_q_net_x0,
    i_15 => delay14_q_net_x0,
    i_16 => delay15_q_net_x0,
    o => concat1_y_net_x1
  );
  vector_to_scalar1 : entity xil_defaultlib.psb3_0_vector_to_scalar1_x3 
  port map (
    i_1 => delay0_q_net,
    i_2 => delay1_q_net,
    i_3 => delay2_q_net,
    i_4 => delay3_q_net,
    i_5 => delay4_q_net,
    i_6 => delay5_q_net,
    i_7 => delay6_q_net,
    i_8 => delay7_q_net,
    i_9 => delay8_q_net,
    i_10 => delay9_q_net,
    i_11 => delay10_q_net,
    i_12 => delay11_q_net,
    i_13 => delay12_q_net,
    i_14 => delay13_q_net,
    i_15 => delay14_q_net,
    i_16 => delay15_q_net,
    o => concat1_y_net_x0
  );
  vector_to_scalar2 : entity xil_defaultlib.psb3_0_vector_to_scalar2_x3 
  port map (
    i_1 => slice0_y_net,
    i_2 => slice1_y_net,
    i_3 => slice2_y_net,
    i_4 => slice3_y_net,
    i_5 => slice4_y_net,
    i_6 => slice5_y_net,
    i_7 => slice6_y_net,
    i_8 => slice7_y_net,
    i_9 => slice8_y_net,
    i_10 => slice9_y_net,
    i_11 => slice10_y_net,
    i_12 => slice11_y_net,
    i_13 => slice12_y_net,
    i_14 => slice13_y_net,
    i_15 => slice14_y_net,
    i_16 => slice15_y_net,
    o => concat1_y_net
  );
  constant17 : entity xil_defaultlib.sysgen_constant_71e89d757c 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant17_op_net
  );
  convert : entity xil_defaultlib.psb3_0_xlconvert 
  generic map (
    bool_conversion => 1,
    din_arith => 1,
    din_bin_pt => 0,
    din_width => 1,
    dout_arith => 1,
    dout_bin_pt => 0,
    dout_width => 1,
    latency => 1,
    overflow => xlWrap,
    quantization => xlTruncate
  )
  port map (
    clr => '0',
    en => "1",
    din => expression_dout_net,
    clk => clk_net,
    ce => ce_net,
    dout => convert_dout_net
  );
  expression : entity xil_defaultlib.sysgen_expr_7c83532765 
  port map (
    clr => '0',
    a => concat1_y_net_x1,
    b => concat1_y_net_x0,
    s => concat1_y_net,
    clk => clk_net,
    ce => ce_net,
    dout => expression_dout_net
  );
  register_x0 : entity xil_defaultlib.psb3_0_xlregister 
  generic map (
    d_width => 1,
    init_value => b"0"
  )
  port map (
    d => constant17_op_net,
    rst => gin_tl_reset_net,
    en => convert_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => register_q_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Overflow Detector add_re_2/Vector Delay
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_delay_x4 is
  port (
    d_1 : in std_logic_vector( 1-1 downto 0 );
    d_2 : in std_logic_vector( 1-1 downto 0 );
    d_3 : in std_logic_vector( 1-1 downto 0 );
    d_4 : in std_logic_vector( 1-1 downto 0 );
    d_5 : in std_logic_vector( 1-1 downto 0 );
    d_6 : in std_logic_vector( 1-1 downto 0 );
    d_7 : in std_logic_vector( 1-1 downto 0 );
    d_8 : in std_logic_vector( 1-1 downto 0 );
    d_9 : in std_logic_vector( 1-1 downto 0 );
    d_10 : in std_logic_vector( 1-1 downto 0 );
    d_11 : in std_logic_vector( 1-1 downto 0 );
    d_12 : in std_logic_vector( 1-1 downto 0 );
    d_13 : in std_logic_vector( 1-1 downto 0 );
    d_14 : in std_logic_vector( 1-1 downto 0 );
    d_15 : in std_logic_vector( 1-1 downto 0 );
    d_16 : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    q_1 : out std_logic_vector( 1-1 downto 0 );
    q_2 : out std_logic_vector( 1-1 downto 0 );
    q_3 : out std_logic_vector( 1-1 downto 0 );
    q_4 : out std_logic_vector( 1-1 downto 0 );
    q_5 : out std_logic_vector( 1-1 downto 0 );
    q_6 : out std_logic_vector( 1-1 downto 0 );
    q_7 : out std_logic_vector( 1-1 downto 0 );
    q_8 : out std_logic_vector( 1-1 downto 0 );
    q_9 : out std_logic_vector( 1-1 downto 0 );
    q_10 : out std_logic_vector( 1-1 downto 0 );
    q_11 : out std_logic_vector( 1-1 downto 0 );
    q_12 : out std_logic_vector( 1-1 downto 0 );
    q_13 : out std_logic_vector( 1-1 downto 0 );
    q_14 : out std_logic_vector( 1-1 downto 0 );
    q_15 : out std_logic_vector( 1-1 downto 0 );
    q_16 : out std_logic_vector( 1-1 downto 0 )
  );
end psb3_0_vector_delay_x4;
architecture structural of psb3_0_vector_delay_x4 is 
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay0_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay12_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal delay5_q_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal delay8_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay11_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay13_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay7_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay10_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay15_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay14_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay9_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 1-1 downto 0 );
begin
  q_1 <= delay0_q_net;
  q_2 <= delay1_q_net;
  q_3 <= delay2_q_net;
  q_4 <= delay3_q_net;
  q_5 <= delay4_q_net;
  q_6 <= delay5_q_net;
  q_7 <= delay6_q_net;
  q_8 <= delay7_q_net;
  q_9 <= delay8_q_net;
  q_10 <= delay9_q_net;
  q_11 <= delay10_q_net;
  q_12 <= delay11_q_net;
  q_13 <= delay12_q_net;
  q_14 <= delay13_q_net;
  q_15 <= delay14_q_net;
  q_16 <= delay15_q_net;
  slice0_y_net <= d_1;
  slice1_y_net <= d_2;
  slice2_y_net <= d_3;
  slice3_y_net <= d_4;
  slice4_y_net <= d_5;
  slice5_y_net <= d_6;
  slice6_y_net <= d_7;
  slice7_y_net <= d_8;
  slice8_y_net <= d_9;
  slice9_y_net <= d_10;
  slice10_y_net <= d_11;
  slice11_y_net <= d_12;
  slice12_y_net <= d_13;
  slice13_y_net <= d_14;
  slice14_y_net <= d_15;
  slice15_y_net <= d_16;
  clk_net <= clk_1;
  ce_net <= ce_1;
  delay0 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice0_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay0_q_net
  );
  delay1 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice2_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay3 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice3_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  delay4 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice4_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net
  );
  delay5 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice5_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  delay6 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice6_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay6_q_net
  );
  delay7 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice7_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay7_q_net
  );
  delay8 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice8_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay8_q_net
  );
  delay9 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice9_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay9_q_net
  );
  delay10 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice10_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay10_q_net
  );
  delay11 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice11_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay11_q_net
  );
  delay12 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice12_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay12_q_net
  );
  delay13 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice13_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay13_q_net
  );
  delay14 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice14_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay14_q_net
  );
  delay15 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice15_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay15_q_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Overflow Detector add_re_2/Vector Delay1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_delay1_x4 is
  port (
    d_1 : in std_logic_vector( 1-1 downto 0 );
    d_2 : in std_logic_vector( 1-1 downto 0 );
    d_3 : in std_logic_vector( 1-1 downto 0 );
    d_4 : in std_logic_vector( 1-1 downto 0 );
    d_5 : in std_logic_vector( 1-1 downto 0 );
    d_6 : in std_logic_vector( 1-1 downto 0 );
    d_7 : in std_logic_vector( 1-1 downto 0 );
    d_8 : in std_logic_vector( 1-1 downto 0 );
    d_9 : in std_logic_vector( 1-1 downto 0 );
    d_10 : in std_logic_vector( 1-1 downto 0 );
    d_11 : in std_logic_vector( 1-1 downto 0 );
    d_12 : in std_logic_vector( 1-1 downto 0 );
    d_13 : in std_logic_vector( 1-1 downto 0 );
    d_14 : in std_logic_vector( 1-1 downto 0 );
    d_15 : in std_logic_vector( 1-1 downto 0 );
    d_16 : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    q_1 : out std_logic_vector( 1-1 downto 0 );
    q_2 : out std_logic_vector( 1-1 downto 0 );
    q_3 : out std_logic_vector( 1-1 downto 0 );
    q_4 : out std_logic_vector( 1-1 downto 0 );
    q_5 : out std_logic_vector( 1-1 downto 0 );
    q_6 : out std_logic_vector( 1-1 downto 0 );
    q_7 : out std_logic_vector( 1-1 downto 0 );
    q_8 : out std_logic_vector( 1-1 downto 0 );
    q_9 : out std_logic_vector( 1-1 downto 0 );
    q_10 : out std_logic_vector( 1-1 downto 0 );
    q_11 : out std_logic_vector( 1-1 downto 0 );
    q_12 : out std_logic_vector( 1-1 downto 0 );
    q_13 : out std_logic_vector( 1-1 downto 0 );
    q_14 : out std_logic_vector( 1-1 downto 0 );
    q_15 : out std_logic_vector( 1-1 downto 0 );
    q_16 : out std_logic_vector( 1-1 downto 0 )
  );
end psb3_0_vector_delay1_x4;
architecture structural of psb3_0_vector_delay1_x4 is 
  signal delay0_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay7_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay14_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay12_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay15_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay13_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay9_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay10_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay11_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal slice7_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal slice8_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 1-1 downto 0 );
begin
  q_1 <= delay0_q_net;
  q_2 <= delay1_q_net;
  q_3 <= delay2_q_net;
  q_4 <= delay3_q_net;
  q_5 <= delay4_q_net;
  q_6 <= delay5_q_net;
  q_7 <= delay6_q_net;
  q_8 <= delay7_q_net;
  q_9 <= delay8_q_net;
  q_10 <= delay9_q_net;
  q_11 <= delay10_q_net;
  q_12 <= delay11_q_net;
  q_13 <= delay12_q_net;
  q_14 <= delay13_q_net;
  q_15 <= delay14_q_net;
  q_16 <= delay15_q_net;
  slice0_y_net <= d_1;
  slice1_y_net <= d_2;
  slice2_y_net <= d_3;
  slice3_y_net <= d_4;
  slice4_y_net <= d_5;
  slice5_y_net <= d_6;
  slice6_y_net <= d_7;
  slice7_y_net <= d_8;
  slice8_y_net <= d_9;
  slice9_y_net <= d_10;
  slice10_y_net <= d_11;
  slice11_y_net <= d_12;
  slice12_y_net <= d_13;
  slice13_y_net <= d_14;
  slice14_y_net <= d_15;
  slice15_y_net <= d_16;
  clk_net <= clk_1;
  ce_net <= ce_1;
  delay0 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice0_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay0_q_net
  );
  delay1 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice2_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay3 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice3_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  delay4 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice4_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net
  );
  delay5 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice5_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  delay6 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice6_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay6_q_net
  );
  delay7 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice7_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay7_q_net
  );
  delay8 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice8_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay8_q_net
  );
  delay9 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice9_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay9_q_net
  );
  delay10 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice10_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay10_q_net
  );
  delay11 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice11_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay11_q_net
  );
  delay12 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice12_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay12_q_net
  );
  delay13 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice13_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay13_q_net
  );
  delay14 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice14_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay14_q_net
  );
  delay15 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice15_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay15_q_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Overflow Detector add_re_2/Vector Slice
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_slice_x4 is
  port (
    in_1 : in std_logic_vector( 16-1 downto 0 );
    in_2 : in std_logic_vector( 16-1 downto 0 );
    in_3 : in std_logic_vector( 16-1 downto 0 );
    in_4 : in std_logic_vector( 16-1 downto 0 );
    in_5 : in std_logic_vector( 16-1 downto 0 );
    in_6 : in std_logic_vector( 16-1 downto 0 );
    in_7 : in std_logic_vector( 16-1 downto 0 );
    in_8 : in std_logic_vector( 16-1 downto 0 );
    in_9 : in std_logic_vector( 16-1 downto 0 );
    in_10 : in std_logic_vector( 16-1 downto 0 );
    in_11 : in std_logic_vector( 16-1 downto 0 );
    in_12 : in std_logic_vector( 16-1 downto 0 );
    in_13 : in std_logic_vector( 16-1 downto 0 );
    in_14 : in std_logic_vector( 16-1 downto 0 );
    in_15 : in std_logic_vector( 16-1 downto 0 );
    in_16 : in std_logic_vector( 16-1 downto 0 );
    out_1 : out std_logic_vector( 1-1 downto 0 );
    out_2 : out std_logic_vector( 1-1 downto 0 );
    out_3 : out std_logic_vector( 1-1 downto 0 );
    out_4 : out std_logic_vector( 1-1 downto 0 );
    out_5 : out std_logic_vector( 1-1 downto 0 );
    out_6 : out std_logic_vector( 1-1 downto 0 );
    out_7 : out std_logic_vector( 1-1 downto 0 );
    out_8 : out std_logic_vector( 1-1 downto 0 );
    out_9 : out std_logic_vector( 1-1 downto 0 );
    out_10 : out std_logic_vector( 1-1 downto 0 );
    out_11 : out std_logic_vector( 1-1 downto 0 );
    out_12 : out std_logic_vector( 1-1 downto 0 );
    out_13 : out std_logic_vector( 1-1 downto 0 );
    out_14 : out std_logic_vector( 1-1 downto 0 );
    out_15 : out std_logic_vector( 1-1 downto 0 );
    out_16 : out std_logic_vector( 1-1 downto 0 )
  );
end psb3_0_vector_slice_x4;
architecture structural of psb3_0_vector_slice_x4 is 
  signal mult13_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult14_p_net : std_logic_vector( 16-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 1-1 downto 0 );
  signal mult3_p_net : std_logic_vector( 16-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 1-1 downto 0 );
  signal mult5_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult8_p_net : std_logic_vector( 16-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 1-1 downto 0 );
  signal mult4_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult6_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult7_p_net : std_logic_vector( 16-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 1-1 downto 0 );
  signal mult1_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult9_p_net : std_logic_vector( 16-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 1-1 downto 0 );
  signal mult2_p_net : std_logic_vector( 16-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 1-1 downto 0 );
  signal mult10_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult0_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult11_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult12_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult15_p_net : std_logic_vector( 16-1 downto 0 );
begin
  out_1 <= slice0_y_net;
  out_2 <= slice1_y_net;
  out_3 <= slice2_y_net;
  out_4 <= slice3_y_net;
  out_5 <= slice4_y_net;
  out_6 <= slice5_y_net;
  out_7 <= slice6_y_net;
  out_8 <= slice7_y_net;
  out_9 <= slice8_y_net;
  out_10 <= slice9_y_net;
  out_11 <= slice10_y_net;
  out_12 <= slice11_y_net;
  out_13 <= slice12_y_net;
  out_14 <= slice13_y_net;
  out_15 <= slice14_y_net;
  out_16 <= slice15_y_net;
  mult0_p_net <= in_1;
  mult1_p_net <= in_2;
  mult2_p_net <= in_3;
  mult3_p_net <= in_4;
  mult4_p_net <= in_5;
  mult5_p_net <= in_6;
  mult6_p_net <= in_7;
  mult7_p_net <= in_8;
  mult8_p_net <= in_9;
  mult9_p_net <= in_10;
  mult10_p_net <= in_11;
  mult11_p_net <= in_12;
  mult12_p_net <= in_13;
  mult13_p_net <= in_14;
  mult14_p_net <= in_15;
  mult15_p_net <= in_16;
  slice0 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult0_p_net,
    y => slice0_y_net
  );
  slice1 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult1_p_net,
    y => slice1_y_net
  );
  slice2 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult2_p_net,
    y => slice2_y_net
  );
  slice3 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult3_p_net,
    y => slice3_y_net
  );
  slice4 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult4_p_net,
    y => slice4_y_net
  );
  slice5 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult5_p_net,
    y => slice5_y_net
  );
  slice6 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult6_p_net,
    y => slice6_y_net
  );
  slice7 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult7_p_net,
    y => slice7_y_net
  );
  slice8 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult8_p_net,
    y => slice8_y_net
  );
  slice9 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult9_p_net,
    y => slice9_y_net
  );
  slice10 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult10_p_net,
    y => slice10_y_net
  );
  slice11 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult11_p_net,
    y => slice11_y_net
  );
  slice12 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult12_p_net,
    y => slice12_y_net
  );
  slice13 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult13_p_net,
    y => slice13_y_net
  );
  slice14 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult14_p_net,
    y => slice14_y_net
  );
  slice15 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult15_p_net,
    y => slice15_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Overflow Detector add_re_2/Vector Slice1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_slice1_x4 is
  port (
    in_1 : in std_logic_vector( 16-1 downto 0 );
    in_2 : in std_logic_vector( 16-1 downto 0 );
    in_3 : in std_logic_vector( 16-1 downto 0 );
    in_4 : in std_logic_vector( 16-1 downto 0 );
    in_5 : in std_logic_vector( 16-1 downto 0 );
    in_6 : in std_logic_vector( 16-1 downto 0 );
    in_7 : in std_logic_vector( 16-1 downto 0 );
    in_8 : in std_logic_vector( 16-1 downto 0 );
    in_9 : in std_logic_vector( 16-1 downto 0 );
    in_10 : in std_logic_vector( 16-1 downto 0 );
    in_11 : in std_logic_vector( 16-1 downto 0 );
    in_12 : in std_logic_vector( 16-1 downto 0 );
    in_13 : in std_logic_vector( 16-1 downto 0 );
    in_14 : in std_logic_vector( 16-1 downto 0 );
    in_15 : in std_logic_vector( 16-1 downto 0 );
    in_16 : in std_logic_vector( 16-1 downto 0 );
    out_1 : out std_logic_vector( 1-1 downto 0 );
    out_2 : out std_logic_vector( 1-1 downto 0 );
    out_3 : out std_logic_vector( 1-1 downto 0 );
    out_4 : out std_logic_vector( 1-1 downto 0 );
    out_5 : out std_logic_vector( 1-1 downto 0 );
    out_6 : out std_logic_vector( 1-1 downto 0 );
    out_7 : out std_logic_vector( 1-1 downto 0 );
    out_8 : out std_logic_vector( 1-1 downto 0 );
    out_9 : out std_logic_vector( 1-1 downto 0 );
    out_10 : out std_logic_vector( 1-1 downto 0 );
    out_11 : out std_logic_vector( 1-1 downto 0 );
    out_12 : out std_logic_vector( 1-1 downto 0 );
    out_13 : out std_logic_vector( 1-1 downto 0 );
    out_14 : out std_logic_vector( 1-1 downto 0 );
    out_15 : out std_logic_vector( 1-1 downto 0 );
    out_16 : out std_logic_vector( 1-1 downto 0 )
  );
end psb3_0_vector_slice1_x4;
architecture structural of psb3_0_vector_slice1_x4 is 
  signal slice1_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
begin
  out_1 <= slice0_y_net;
  out_2 <= slice1_y_net;
  out_3 <= slice2_y_net;
  out_4 <= slice3_y_net;
  out_5 <= slice4_y_net;
  out_6 <= slice5_y_net;
  out_7 <= slice6_y_net;
  out_8 <= slice7_y_net;
  out_9 <= slice8_y_net;
  out_10 <= slice9_y_net;
  out_11 <= slice10_y_net;
  out_12 <= slice11_y_net;
  out_13 <= slice12_y_net;
  out_14 <= slice13_y_net;
  out_15 <= slice14_y_net;
  out_16 <= slice15_y_net;
  reinterpret0_output_port_net <= in_1;
  reinterpret1_output_port_net <= in_2;
  reinterpret2_output_port_net <= in_3;
  reinterpret3_output_port_net <= in_4;
  reinterpret4_output_port_net <= in_5;
  reinterpret5_output_port_net <= in_6;
  reinterpret6_output_port_net <= in_7;
  reinterpret7_output_port_net <= in_8;
  reinterpret8_output_port_net <= in_9;
  reinterpret9_output_port_net <= in_10;
  reinterpret10_output_port_net <= in_11;
  reinterpret11_output_port_net <= in_12;
  reinterpret12_output_port_net <= in_13;
  reinterpret13_output_port_net <= in_14;
  reinterpret14_output_port_net <= in_15;
  reinterpret15_output_port_net <= in_16;
  slice0 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret0_output_port_net,
    y => slice0_y_net
  );
  slice1 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret1_output_port_net,
    y => slice1_y_net
  );
  slice2 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret2_output_port_net,
    y => slice2_y_net
  );
  slice3 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret3_output_port_net,
    y => slice3_y_net
  );
  slice4 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret4_output_port_net,
    y => slice4_y_net
  );
  slice5 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret5_output_port_net,
    y => slice5_y_net
  );
  slice6 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret6_output_port_net,
    y => slice6_y_net
  );
  slice7 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret7_output_port_net,
    y => slice7_y_net
  );
  slice8 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret8_output_port_net,
    y => slice8_y_net
  );
  slice9 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret9_output_port_net,
    y => slice9_y_net
  );
  slice10 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret10_output_port_net,
    y => slice10_y_net
  );
  slice11 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret11_output_port_net,
    y => slice11_y_net
  );
  slice12 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret12_output_port_net,
    y => slice12_y_net
  );
  slice13 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret13_output_port_net,
    y => slice13_y_net
  );
  slice14 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret14_output_port_net,
    y => slice14_y_net
  );
  slice15 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret15_output_port_net,
    y => slice15_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Overflow Detector add_re_2/Vector Slice2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_slice2_x4 is
  port (
    in_1 : in std_logic_vector( 16-1 downto 0 );
    in_2 : in std_logic_vector( 16-1 downto 0 );
    in_3 : in std_logic_vector( 16-1 downto 0 );
    in_4 : in std_logic_vector( 16-1 downto 0 );
    in_5 : in std_logic_vector( 16-1 downto 0 );
    in_6 : in std_logic_vector( 16-1 downto 0 );
    in_7 : in std_logic_vector( 16-1 downto 0 );
    in_8 : in std_logic_vector( 16-1 downto 0 );
    in_9 : in std_logic_vector( 16-1 downto 0 );
    in_10 : in std_logic_vector( 16-1 downto 0 );
    in_11 : in std_logic_vector( 16-1 downto 0 );
    in_12 : in std_logic_vector( 16-1 downto 0 );
    in_13 : in std_logic_vector( 16-1 downto 0 );
    in_14 : in std_logic_vector( 16-1 downto 0 );
    in_15 : in std_logic_vector( 16-1 downto 0 );
    in_16 : in std_logic_vector( 16-1 downto 0 );
    out_1 : out std_logic_vector( 1-1 downto 0 );
    out_2 : out std_logic_vector( 1-1 downto 0 );
    out_3 : out std_logic_vector( 1-1 downto 0 );
    out_4 : out std_logic_vector( 1-1 downto 0 );
    out_5 : out std_logic_vector( 1-1 downto 0 );
    out_6 : out std_logic_vector( 1-1 downto 0 );
    out_7 : out std_logic_vector( 1-1 downto 0 );
    out_8 : out std_logic_vector( 1-1 downto 0 );
    out_9 : out std_logic_vector( 1-1 downto 0 );
    out_10 : out std_logic_vector( 1-1 downto 0 );
    out_11 : out std_logic_vector( 1-1 downto 0 );
    out_12 : out std_logic_vector( 1-1 downto 0 );
    out_13 : out std_logic_vector( 1-1 downto 0 );
    out_14 : out std_logic_vector( 1-1 downto 0 );
    out_15 : out std_logic_vector( 1-1 downto 0 );
    out_16 : out std_logic_vector( 1-1 downto 0 )
  );
end psb3_0_vector_slice2_x4;
architecture structural of psb3_0_vector_slice2_x4 is 
  signal addsub2_s_net : std_logic_vector( 16-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 1-1 downto 0 );
  signal addsub8_s_net : std_logic_vector( 16-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 1-1 downto 0 );
  signal addsub10_s_net : std_logic_vector( 16-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 1-1 downto 0 );
  signal addsub11_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub13_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub6_s_net : std_logic_vector( 16-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 1-1 downto 0 );
  signal addsub5_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub12_s_net : std_logic_vector( 16-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 1-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 16-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 1-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 16-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 1-1 downto 0 );
  signal addsub7_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub3_s_net : std_logic_vector( 16-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 1-1 downto 0 );
  signal addsub9_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub0_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub15_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub14_s_net : std_logic_vector( 16-1 downto 0 );
begin
  out_1 <= slice0_y_net;
  out_2 <= slice1_y_net;
  out_3 <= slice2_y_net;
  out_4 <= slice3_y_net;
  out_5 <= slice4_y_net;
  out_6 <= slice5_y_net;
  out_7 <= slice6_y_net;
  out_8 <= slice7_y_net;
  out_9 <= slice8_y_net;
  out_10 <= slice9_y_net;
  out_11 <= slice10_y_net;
  out_12 <= slice11_y_net;
  out_13 <= slice12_y_net;
  out_14 <= slice13_y_net;
  out_15 <= slice14_y_net;
  out_16 <= slice15_y_net;
  addsub0_s_net <= in_1;
  addsub1_s_net <= in_2;
  addsub2_s_net <= in_3;
  addsub3_s_net <= in_4;
  addsub4_s_net <= in_5;
  addsub5_s_net <= in_6;
  addsub6_s_net <= in_7;
  addsub7_s_net <= in_8;
  addsub8_s_net <= in_9;
  addsub9_s_net <= in_10;
  addsub10_s_net <= in_11;
  addsub11_s_net <= in_12;
  addsub12_s_net <= in_13;
  addsub13_s_net <= in_14;
  addsub14_s_net <= in_15;
  addsub15_s_net <= in_16;
  slice0 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub0_s_net,
    y => slice0_y_net
  );
  slice1 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub1_s_net,
    y => slice1_y_net
  );
  slice2 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub2_s_net,
    y => slice2_y_net
  );
  slice3 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub3_s_net,
    y => slice3_y_net
  );
  slice4 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub4_s_net,
    y => slice4_y_net
  );
  slice5 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub5_s_net,
    y => slice5_y_net
  );
  slice6 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub6_s_net,
    y => slice6_y_net
  );
  slice7 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub7_s_net,
    y => slice7_y_net
  );
  slice8 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub8_s_net,
    y => slice8_y_net
  );
  slice9 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub9_s_net,
    y => slice9_y_net
  );
  slice10 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub10_s_net,
    y => slice10_y_net
  );
  slice11 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub11_s_net,
    y => slice11_y_net
  );
  slice12 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub12_s_net,
    y => slice12_y_net
  );
  slice13 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub13_s_net,
    y => slice13_y_net
  );
  slice14 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub14_s_net,
    y => slice14_y_net
  );
  slice15 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub15_s_net,
    y => slice15_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Overflow Detector add_re_2/Vector to Scalar
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_to_scalar_x4 is
  port (
    i_1 : in std_logic_vector( 1-1 downto 0 );
    i_2 : in std_logic_vector( 1-1 downto 0 );
    i_3 : in std_logic_vector( 1-1 downto 0 );
    i_4 : in std_logic_vector( 1-1 downto 0 );
    i_5 : in std_logic_vector( 1-1 downto 0 );
    i_6 : in std_logic_vector( 1-1 downto 0 );
    i_7 : in std_logic_vector( 1-1 downto 0 );
    i_8 : in std_logic_vector( 1-1 downto 0 );
    i_9 : in std_logic_vector( 1-1 downto 0 );
    i_10 : in std_logic_vector( 1-1 downto 0 );
    i_11 : in std_logic_vector( 1-1 downto 0 );
    i_12 : in std_logic_vector( 1-1 downto 0 );
    i_13 : in std_logic_vector( 1-1 downto 0 );
    i_14 : in std_logic_vector( 1-1 downto 0 );
    i_15 : in std_logic_vector( 1-1 downto 0 );
    i_16 : in std_logic_vector( 1-1 downto 0 );
    o : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_vector_to_scalar_x4;
architecture structural of psb3_0_vector_to_scalar_x4 is 
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay7_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 1-1 downto 0 );
  signal concat1_y_net : std_logic_vector( 16-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay9_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay11_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay10_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay12_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay0_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay15_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay14_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay13_q_net : std_logic_vector( 1-1 downto 0 );
begin
  o <= concat1_y_net;
  delay0_q_net <= i_1;
  delay1_q_net <= i_2;
  delay2_q_net <= i_3;
  delay3_q_net <= i_4;
  delay4_q_net <= i_5;
  delay5_q_net <= i_6;
  delay6_q_net <= i_7;
  delay7_q_net <= i_8;
  delay8_q_net <= i_9;
  delay9_q_net <= i_10;
  delay10_q_net <= i_11;
  delay11_q_net <= i_12;
  delay12_q_net <= i_13;
  delay13_q_net <= i_14;
  delay14_q_net <= i_15;
  delay15_q_net <= i_16;
  concat1 : entity xil_defaultlib.sysgen_concat_d977c66e35 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => delay15_q_net,
    in1 => delay14_q_net,
    in2 => delay13_q_net,
    in3 => delay12_q_net,
    in4 => delay11_q_net,
    in5 => delay10_q_net,
    in6 => delay9_q_net,
    in7 => delay8_q_net,
    in8 => delay7_q_net,
    in9 => delay6_q_net,
    in10 => delay5_q_net,
    in11 => delay4_q_net,
    in12 => delay3_q_net,
    in13 => delay2_q_net,
    in14 => delay1_q_net,
    in15 => delay0_q_net,
    y => concat1_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Overflow Detector add_re_2/Vector to Scalar1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_to_scalar1_x4 is
  port (
    i_1 : in std_logic_vector( 1-1 downto 0 );
    i_2 : in std_logic_vector( 1-1 downto 0 );
    i_3 : in std_logic_vector( 1-1 downto 0 );
    i_4 : in std_logic_vector( 1-1 downto 0 );
    i_5 : in std_logic_vector( 1-1 downto 0 );
    i_6 : in std_logic_vector( 1-1 downto 0 );
    i_7 : in std_logic_vector( 1-1 downto 0 );
    i_8 : in std_logic_vector( 1-1 downto 0 );
    i_9 : in std_logic_vector( 1-1 downto 0 );
    i_10 : in std_logic_vector( 1-1 downto 0 );
    i_11 : in std_logic_vector( 1-1 downto 0 );
    i_12 : in std_logic_vector( 1-1 downto 0 );
    i_13 : in std_logic_vector( 1-1 downto 0 );
    i_14 : in std_logic_vector( 1-1 downto 0 );
    i_15 : in std_logic_vector( 1-1 downto 0 );
    i_16 : in std_logic_vector( 1-1 downto 0 );
    o : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_vector_to_scalar1_x4;
architecture structural of psb3_0_vector_to_scalar1_x4 is 
  signal delay0_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay12_q_net : std_logic_vector( 1-1 downto 0 );
  signal concat1_y_net : std_logic_vector( 16-1 downto 0 );
  signal delay14_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay15_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay11_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay10_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay13_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay9_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay7_q_net : std_logic_vector( 1-1 downto 0 );
begin
  o <= concat1_y_net;
  delay0_q_net <= i_1;
  delay1_q_net <= i_2;
  delay2_q_net <= i_3;
  delay3_q_net <= i_4;
  delay4_q_net <= i_5;
  delay5_q_net <= i_6;
  delay6_q_net <= i_7;
  delay7_q_net <= i_8;
  delay8_q_net <= i_9;
  delay9_q_net <= i_10;
  delay10_q_net <= i_11;
  delay11_q_net <= i_12;
  delay12_q_net <= i_13;
  delay13_q_net <= i_14;
  delay14_q_net <= i_15;
  delay15_q_net <= i_16;
  concat1 : entity xil_defaultlib.sysgen_concat_d977c66e35 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => delay15_q_net,
    in1 => delay14_q_net,
    in2 => delay13_q_net,
    in3 => delay12_q_net,
    in4 => delay11_q_net,
    in5 => delay10_q_net,
    in6 => delay9_q_net,
    in7 => delay8_q_net,
    in8 => delay7_q_net,
    in9 => delay6_q_net,
    in10 => delay5_q_net,
    in11 => delay4_q_net,
    in12 => delay3_q_net,
    in13 => delay2_q_net,
    in14 => delay1_q_net,
    in15 => delay0_q_net,
    y => concat1_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Overflow Detector add_re_2/Vector to Scalar2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_to_scalar2_x4 is
  port (
    i_1 : in std_logic_vector( 1-1 downto 0 );
    i_2 : in std_logic_vector( 1-1 downto 0 );
    i_3 : in std_logic_vector( 1-1 downto 0 );
    i_4 : in std_logic_vector( 1-1 downto 0 );
    i_5 : in std_logic_vector( 1-1 downto 0 );
    i_6 : in std_logic_vector( 1-1 downto 0 );
    i_7 : in std_logic_vector( 1-1 downto 0 );
    i_8 : in std_logic_vector( 1-1 downto 0 );
    i_9 : in std_logic_vector( 1-1 downto 0 );
    i_10 : in std_logic_vector( 1-1 downto 0 );
    i_11 : in std_logic_vector( 1-1 downto 0 );
    i_12 : in std_logic_vector( 1-1 downto 0 );
    i_13 : in std_logic_vector( 1-1 downto 0 );
    i_14 : in std_logic_vector( 1-1 downto 0 );
    i_15 : in std_logic_vector( 1-1 downto 0 );
    i_16 : in std_logic_vector( 1-1 downto 0 );
    o : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_vector_to_scalar2_x4;
architecture structural of psb3_0_vector_to_scalar2_x4 is 
  signal slice6_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 1-1 downto 0 );
  signal concat1_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 1-1 downto 0 );
begin
  o <= concat1_y_net;
  slice0_y_net <= i_1;
  slice1_y_net <= i_2;
  slice2_y_net <= i_3;
  slice3_y_net <= i_4;
  slice4_y_net <= i_5;
  slice5_y_net <= i_6;
  slice6_y_net <= i_7;
  slice7_y_net <= i_8;
  slice8_y_net <= i_9;
  slice9_y_net <= i_10;
  slice10_y_net <= i_11;
  slice11_y_net <= i_12;
  slice12_y_net <= i_13;
  slice13_y_net <= i_14;
  slice14_y_net <= i_15;
  slice15_y_net <= i_16;
  concat1 : entity xil_defaultlib.sysgen_concat_d977c66e35 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => slice15_y_net,
    in1 => slice14_y_net,
    in2 => slice13_y_net,
    in3 => slice12_y_net,
    in4 => slice11_y_net,
    in5 => slice10_y_net,
    in6 => slice9_y_net,
    in7 => slice8_y_net,
    in8 => slice7_y_net,
    in9 => slice6_y_net,
    in10 => slice5_y_net,
    in11 => slice4_y_net,
    in12 => slice3_y_net,
    in13 => slice2_y_net,
    in14 => slice1_y_net,
    in15 => slice0_y_net,
    y => concat1_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Overflow Detector add_re_2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_overflow_detector_add_re_2 is
  port (
    rst : in std_logic_vector( 1-1 downto 0 );
    a_1 : in std_logic_vector( 16-1 downto 0 );
    b_1 : in std_logic_vector( 16-1 downto 0 );
    s_1 : in std_logic_vector( 16-1 downto 0 );
    a_2 : in std_logic_vector( 16-1 downto 0 );
    a_3 : in std_logic_vector( 16-1 downto 0 );
    a_4 : in std_logic_vector( 16-1 downto 0 );
    a_5 : in std_logic_vector( 16-1 downto 0 );
    a_6 : in std_logic_vector( 16-1 downto 0 );
    a_7 : in std_logic_vector( 16-1 downto 0 );
    a_8 : in std_logic_vector( 16-1 downto 0 );
    a_9 : in std_logic_vector( 16-1 downto 0 );
    a_10 : in std_logic_vector( 16-1 downto 0 );
    a_11 : in std_logic_vector( 16-1 downto 0 );
    a_12 : in std_logic_vector( 16-1 downto 0 );
    a_13 : in std_logic_vector( 16-1 downto 0 );
    a_14 : in std_logic_vector( 16-1 downto 0 );
    a_15 : in std_logic_vector( 16-1 downto 0 );
    a_16 : in std_logic_vector( 16-1 downto 0 );
    b_2 : in std_logic_vector( 16-1 downto 0 );
    b_3 : in std_logic_vector( 16-1 downto 0 );
    b_4 : in std_logic_vector( 16-1 downto 0 );
    b_5 : in std_logic_vector( 16-1 downto 0 );
    b_6 : in std_logic_vector( 16-1 downto 0 );
    b_7 : in std_logic_vector( 16-1 downto 0 );
    b_8 : in std_logic_vector( 16-1 downto 0 );
    b_9 : in std_logic_vector( 16-1 downto 0 );
    b_10 : in std_logic_vector( 16-1 downto 0 );
    b_11 : in std_logic_vector( 16-1 downto 0 );
    b_12 : in std_logic_vector( 16-1 downto 0 );
    b_13 : in std_logic_vector( 16-1 downto 0 );
    b_14 : in std_logic_vector( 16-1 downto 0 );
    b_15 : in std_logic_vector( 16-1 downto 0 );
    b_16 : in std_logic_vector( 16-1 downto 0 );
    s_2 : in std_logic_vector( 16-1 downto 0 );
    s_3 : in std_logic_vector( 16-1 downto 0 );
    s_4 : in std_logic_vector( 16-1 downto 0 );
    s_5 : in std_logic_vector( 16-1 downto 0 );
    s_6 : in std_logic_vector( 16-1 downto 0 );
    s_7 : in std_logic_vector( 16-1 downto 0 );
    s_8 : in std_logic_vector( 16-1 downto 0 );
    s_9 : in std_logic_vector( 16-1 downto 0 );
    s_10 : in std_logic_vector( 16-1 downto 0 );
    s_11 : in std_logic_vector( 16-1 downto 0 );
    s_12 : in std_logic_vector( 16-1 downto 0 );
    s_13 : in std_logic_vector( 16-1 downto 0 );
    s_14 : in std_logic_vector( 16-1 downto 0 );
    s_15 : in std_logic_vector( 16-1 downto 0 );
    s_16 : in std_logic_vector( 16-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    ov : out std_logic_vector( 1-1 downto 0 )
  );
end psb3_0_overflow_detector_add_re_2;
architecture structural of psb3_0_overflow_detector_add_re_2 is 
  signal mult1_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult10_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mult5_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mult9_p_net : std_logic_vector( 16-1 downto 0 );
  signal register_q_net : std_logic_vector( 1-1 downto 0 );
  signal mult4_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult11_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub0_s_net : std_logic_vector( 16-1 downto 0 );
  signal mult2_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult3_p_net : std_logic_vector( 16-1 downto 0 );
  signal gin_tl_reset_net : std_logic_vector( 1-1 downto 0 );
  signal mult13_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult14_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mult6_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult7_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult8_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult0_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult12_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult15_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub15_s_net : std_logic_vector( 16-1 downto 0 );
  signal delay1_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal addsub8_s_net : std_logic_vector( 16-1 downto 0 );
  signal delay4_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay5_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay6_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay11_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal addsub5_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub6_s_net : std_logic_vector( 16-1 downto 0 );
  signal delay12_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay10_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub13_s_net : std_logic_vector( 16-1 downto 0 );
  signal ce_net : std_logic;
  signal delay9_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay14_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal addsub14_s_net : std_logic_vector( 16-1 downto 0 );
  signal delay13_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub3_s_net : std_logic_vector( 16-1 downto 0 );
  signal delay3_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay0_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal addsub11_s_net : std_logic_vector( 16-1 downto 0 );
  signal delay7_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay8_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal addsub10_s_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub12_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub7_s_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal clk_net : std_logic;
  signal delay2_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal addsub9_s_net : std_logic_vector( 16-1 downto 0 );
  signal slice9_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice13_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice5_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal slice10_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay13_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice0_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice4_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice1_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal slice14_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal slice15_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay7_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice14_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice2_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal slice0_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal slice12_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal slice3_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay14_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice1_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice12_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice7_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice2_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice6_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice11_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal slice6_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay12_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice8_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice10_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice15_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice5_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay15_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay15_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice7_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal slice8_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal slice13_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal delay9_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay10_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay0_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay11_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice3_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice11_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice9_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice4_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 1-1 downto 0 );
  signal expression_dout_net : std_logic_vector( 1-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 1-1 downto 0 );
  signal concat1_y_net_x1 : std_logic_vector( 16-1 downto 0 );
  signal convert_dout_net : std_logic_vector( 1-1 downto 0 );
  signal concat1_y_net : std_logic_vector( 16-1 downto 0 );
  signal constant17_op_net : std_logic_vector( 1-1 downto 0 );
  signal concat1_y_net_x0 : std_logic_vector( 16-1 downto 0 );
begin
  ov <= register_q_net;
  gin_tl_reset_net <= rst;
  mult0_p_net <= a_1;
  reinterpret0_output_port_net <= b_1;
  addsub0_s_net <= s_1;
  mult1_p_net <= a_2;
  mult2_p_net <= a_3;
  mult3_p_net <= a_4;
  mult4_p_net <= a_5;
  mult5_p_net <= a_6;
  mult6_p_net <= a_7;
  mult7_p_net <= a_8;
  mult8_p_net <= a_9;
  mult9_p_net <= a_10;
  mult10_p_net <= a_11;
  mult11_p_net <= a_12;
  mult12_p_net <= a_13;
  mult13_p_net <= a_14;
  mult14_p_net <= a_15;
  mult15_p_net <= a_16;
  reinterpret1_output_port_net <= b_2;
  reinterpret2_output_port_net <= b_3;
  reinterpret3_output_port_net <= b_4;
  reinterpret4_output_port_net <= b_5;
  reinterpret5_output_port_net <= b_6;
  reinterpret6_output_port_net <= b_7;
  reinterpret7_output_port_net <= b_8;
  reinterpret8_output_port_net <= b_9;
  reinterpret9_output_port_net <= b_10;
  reinterpret10_output_port_net <= b_11;
  reinterpret11_output_port_net <= b_12;
  reinterpret12_output_port_net <= b_13;
  reinterpret13_output_port_net <= b_14;
  reinterpret14_output_port_net <= b_15;
  reinterpret15_output_port_net <= b_16;
  addsub1_s_net <= s_2;
  addsub2_s_net <= s_3;
  addsub3_s_net <= s_4;
  addsub4_s_net <= s_5;
  addsub5_s_net <= s_6;
  addsub6_s_net <= s_7;
  addsub7_s_net <= s_8;
  addsub8_s_net <= s_9;
  addsub9_s_net <= s_10;
  addsub10_s_net <= s_11;
  addsub11_s_net <= s_12;
  addsub12_s_net <= s_13;
  addsub13_s_net <= s_14;
  addsub14_s_net <= s_15;
  addsub15_s_net <= s_16;
  clk_net <= clk_1;
  ce_net <= ce_1;
  vector_delay : entity xil_defaultlib.psb3_0_vector_delay_x4 
  port map (
    d_1 => slice0_y_net_x1,
    d_2 => slice1_y_net_x1,
    d_3 => slice2_y_net_x1,
    d_4 => slice3_y_net_x1,
    d_5 => slice4_y_net_x1,
    d_6 => slice5_y_net_x1,
    d_7 => slice6_y_net_x1,
    d_8 => slice7_y_net_x1,
    d_9 => slice8_y_net_x1,
    d_10 => slice9_y_net_x1,
    d_11 => slice10_y_net_x1,
    d_12 => slice11_y_net_x1,
    d_13 => slice12_y_net_x1,
    d_14 => slice13_y_net_x1,
    d_15 => slice14_y_net_x1,
    d_16 => slice15_y_net_x1,
    clk_1 => clk_net,
    ce_1 => ce_net,
    q_1 => delay0_q_net_x0,
    q_2 => delay1_q_net_x0,
    q_3 => delay2_q_net_x0,
    q_4 => delay3_q_net_x0,
    q_5 => delay4_q_net_x0,
    q_6 => delay5_q_net_x0,
    q_7 => delay6_q_net_x0,
    q_8 => delay7_q_net_x0,
    q_9 => delay8_q_net_x0,
    q_10 => delay9_q_net_x0,
    q_11 => delay10_q_net_x0,
    q_12 => delay11_q_net_x0,
    q_13 => delay12_q_net_x0,
    q_14 => delay13_q_net_x0,
    q_15 => delay14_q_net_x0,
    q_16 => delay15_q_net_x0
  );
  vector_delay1 : entity xil_defaultlib.psb3_0_vector_delay1_x4 
  port map (
    d_1 => slice0_y_net_x0,
    d_2 => slice1_y_net_x0,
    d_3 => slice2_y_net_x0,
    d_4 => slice3_y_net_x0,
    d_5 => slice4_y_net_x0,
    d_6 => slice5_y_net_x0,
    d_7 => slice6_y_net_x0,
    d_8 => slice7_y_net_x0,
    d_9 => slice8_y_net_x0,
    d_10 => slice9_y_net_x0,
    d_11 => slice10_y_net_x0,
    d_12 => slice11_y_net_x0,
    d_13 => slice12_y_net_x0,
    d_14 => slice13_y_net_x0,
    d_15 => slice14_y_net_x0,
    d_16 => slice15_y_net_x0,
    clk_1 => clk_net,
    ce_1 => ce_net,
    q_1 => delay0_q_net,
    q_2 => delay1_q_net,
    q_3 => delay2_q_net,
    q_4 => delay3_q_net,
    q_5 => delay4_q_net,
    q_6 => delay5_q_net,
    q_7 => delay6_q_net,
    q_8 => delay7_q_net,
    q_9 => delay8_q_net,
    q_10 => delay9_q_net,
    q_11 => delay10_q_net,
    q_12 => delay11_q_net,
    q_13 => delay12_q_net,
    q_14 => delay13_q_net,
    q_15 => delay14_q_net,
    q_16 => delay15_q_net
  );
  vector_slice : entity xil_defaultlib.psb3_0_vector_slice_x4 
  port map (
    in_1 => mult0_p_net,
    in_2 => mult1_p_net,
    in_3 => mult2_p_net,
    in_4 => mult3_p_net,
    in_5 => mult4_p_net,
    in_6 => mult5_p_net,
    in_7 => mult6_p_net,
    in_8 => mult7_p_net,
    in_9 => mult8_p_net,
    in_10 => mult9_p_net,
    in_11 => mult10_p_net,
    in_12 => mult11_p_net,
    in_13 => mult12_p_net,
    in_14 => mult13_p_net,
    in_15 => mult14_p_net,
    in_16 => mult15_p_net,
    out_1 => slice0_y_net_x1,
    out_2 => slice1_y_net_x1,
    out_3 => slice2_y_net_x1,
    out_4 => slice3_y_net_x1,
    out_5 => slice4_y_net_x1,
    out_6 => slice5_y_net_x1,
    out_7 => slice6_y_net_x1,
    out_8 => slice7_y_net_x1,
    out_9 => slice8_y_net_x1,
    out_10 => slice9_y_net_x1,
    out_11 => slice10_y_net_x1,
    out_12 => slice11_y_net_x1,
    out_13 => slice12_y_net_x1,
    out_14 => slice13_y_net_x1,
    out_15 => slice14_y_net_x1,
    out_16 => slice15_y_net_x1
  );
  vector_slice1 : entity xil_defaultlib.psb3_0_vector_slice1_x4 
  port map (
    in_1 => reinterpret0_output_port_net,
    in_2 => reinterpret1_output_port_net,
    in_3 => reinterpret2_output_port_net,
    in_4 => reinterpret3_output_port_net,
    in_5 => reinterpret4_output_port_net,
    in_6 => reinterpret5_output_port_net,
    in_7 => reinterpret6_output_port_net,
    in_8 => reinterpret7_output_port_net,
    in_9 => reinterpret8_output_port_net,
    in_10 => reinterpret9_output_port_net,
    in_11 => reinterpret10_output_port_net,
    in_12 => reinterpret11_output_port_net,
    in_13 => reinterpret12_output_port_net,
    in_14 => reinterpret13_output_port_net,
    in_15 => reinterpret14_output_port_net,
    in_16 => reinterpret15_output_port_net,
    out_1 => slice0_y_net_x0,
    out_2 => slice1_y_net_x0,
    out_3 => slice2_y_net_x0,
    out_4 => slice3_y_net_x0,
    out_5 => slice4_y_net_x0,
    out_6 => slice5_y_net_x0,
    out_7 => slice6_y_net_x0,
    out_8 => slice7_y_net_x0,
    out_9 => slice8_y_net_x0,
    out_10 => slice9_y_net_x0,
    out_11 => slice10_y_net_x0,
    out_12 => slice11_y_net_x0,
    out_13 => slice12_y_net_x0,
    out_14 => slice13_y_net_x0,
    out_15 => slice14_y_net_x0,
    out_16 => slice15_y_net_x0
  );
  vector_slice2 : entity xil_defaultlib.psb3_0_vector_slice2_x4 
  port map (
    in_1 => addsub0_s_net,
    in_2 => addsub1_s_net,
    in_3 => addsub2_s_net,
    in_4 => addsub3_s_net,
    in_5 => addsub4_s_net,
    in_6 => addsub5_s_net,
    in_7 => addsub6_s_net,
    in_8 => addsub7_s_net,
    in_9 => addsub8_s_net,
    in_10 => addsub9_s_net,
    in_11 => addsub10_s_net,
    in_12 => addsub11_s_net,
    in_13 => addsub12_s_net,
    in_14 => addsub13_s_net,
    in_15 => addsub14_s_net,
    in_16 => addsub15_s_net,
    out_1 => slice0_y_net,
    out_2 => slice1_y_net,
    out_3 => slice2_y_net,
    out_4 => slice3_y_net,
    out_5 => slice4_y_net,
    out_6 => slice5_y_net,
    out_7 => slice6_y_net,
    out_8 => slice7_y_net,
    out_9 => slice8_y_net,
    out_10 => slice9_y_net,
    out_11 => slice10_y_net,
    out_12 => slice11_y_net,
    out_13 => slice12_y_net,
    out_14 => slice13_y_net,
    out_15 => slice14_y_net,
    out_16 => slice15_y_net
  );
  vector_to_scalar : entity xil_defaultlib.psb3_0_vector_to_scalar_x4 
  port map (
    i_1 => delay0_q_net_x0,
    i_2 => delay1_q_net_x0,
    i_3 => delay2_q_net_x0,
    i_4 => delay3_q_net_x0,
    i_5 => delay4_q_net_x0,
    i_6 => delay5_q_net_x0,
    i_7 => delay6_q_net_x0,
    i_8 => delay7_q_net_x0,
    i_9 => delay8_q_net_x0,
    i_10 => delay9_q_net_x0,
    i_11 => delay10_q_net_x0,
    i_12 => delay11_q_net_x0,
    i_13 => delay12_q_net_x0,
    i_14 => delay13_q_net_x0,
    i_15 => delay14_q_net_x0,
    i_16 => delay15_q_net_x0,
    o => concat1_y_net_x1
  );
  vector_to_scalar1 : entity xil_defaultlib.psb3_0_vector_to_scalar1_x4 
  port map (
    i_1 => delay0_q_net,
    i_2 => delay1_q_net,
    i_3 => delay2_q_net,
    i_4 => delay3_q_net,
    i_5 => delay4_q_net,
    i_6 => delay5_q_net,
    i_7 => delay6_q_net,
    i_8 => delay7_q_net,
    i_9 => delay8_q_net,
    i_10 => delay9_q_net,
    i_11 => delay10_q_net,
    i_12 => delay11_q_net,
    i_13 => delay12_q_net,
    i_14 => delay13_q_net,
    i_15 => delay14_q_net,
    i_16 => delay15_q_net,
    o => concat1_y_net_x0
  );
  vector_to_scalar2 : entity xil_defaultlib.psb3_0_vector_to_scalar2_x4 
  port map (
    i_1 => slice0_y_net,
    i_2 => slice1_y_net,
    i_3 => slice2_y_net,
    i_4 => slice3_y_net,
    i_5 => slice4_y_net,
    i_6 => slice5_y_net,
    i_7 => slice6_y_net,
    i_8 => slice7_y_net,
    i_9 => slice8_y_net,
    i_10 => slice9_y_net,
    i_11 => slice10_y_net,
    i_12 => slice11_y_net,
    i_13 => slice12_y_net,
    i_14 => slice13_y_net,
    i_15 => slice14_y_net,
    i_16 => slice15_y_net,
    o => concat1_y_net
  );
  constant17 : entity xil_defaultlib.sysgen_constant_71e89d757c 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant17_op_net
  );
  convert : entity xil_defaultlib.psb3_0_xlconvert 
  generic map (
    bool_conversion => 1,
    din_arith => 1,
    din_bin_pt => 0,
    din_width => 1,
    dout_arith => 1,
    dout_bin_pt => 0,
    dout_width => 1,
    latency => 1,
    overflow => xlWrap,
    quantization => xlTruncate
  )
  port map (
    clr => '0',
    en => "1",
    din => expression_dout_net,
    clk => clk_net,
    ce => ce_net,
    dout => convert_dout_net
  );
  expression : entity xil_defaultlib.sysgen_expr_7c83532765 
  port map (
    clr => '0',
    a => concat1_y_net_x1,
    b => concat1_y_net_x0,
    s => concat1_y_net,
    clk => clk_net,
    ce => ce_net,
    dout => expression_dout_net
  );
  register_x0 : entity xil_defaultlib.psb3_0_xlregister 
  generic map (
    d_width => 1,
    init_value => b"0"
  )
  port map (
    d => constant17_op_net,
    rst => gin_tl_reset_net,
    en => convert_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => register_q_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Overflow Detector add_re_3/Vector Delay
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_delay_x5 is
  port (
    d_1 : in std_logic_vector( 1-1 downto 0 );
    d_2 : in std_logic_vector( 1-1 downto 0 );
    d_3 : in std_logic_vector( 1-1 downto 0 );
    d_4 : in std_logic_vector( 1-1 downto 0 );
    d_5 : in std_logic_vector( 1-1 downto 0 );
    d_6 : in std_logic_vector( 1-1 downto 0 );
    d_7 : in std_logic_vector( 1-1 downto 0 );
    d_8 : in std_logic_vector( 1-1 downto 0 );
    d_9 : in std_logic_vector( 1-1 downto 0 );
    d_10 : in std_logic_vector( 1-1 downto 0 );
    d_11 : in std_logic_vector( 1-1 downto 0 );
    d_12 : in std_logic_vector( 1-1 downto 0 );
    d_13 : in std_logic_vector( 1-1 downto 0 );
    d_14 : in std_logic_vector( 1-1 downto 0 );
    d_15 : in std_logic_vector( 1-1 downto 0 );
    d_16 : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    q_1 : out std_logic_vector( 1-1 downto 0 );
    q_2 : out std_logic_vector( 1-1 downto 0 );
    q_3 : out std_logic_vector( 1-1 downto 0 );
    q_4 : out std_logic_vector( 1-1 downto 0 );
    q_5 : out std_logic_vector( 1-1 downto 0 );
    q_6 : out std_logic_vector( 1-1 downto 0 );
    q_7 : out std_logic_vector( 1-1 downto 0 );
    q_8 : out std_logic_vector( 1-1 downto 0 );
    q_9 : out std_logic_vector( 1-1 downto 0 );
    q_10 : out std_logic_vector( 1-1 downto 0 );
    q_11 : out std_logic_vector( 1-1 downto 0 );
    q_12 : out std_logic_vector( 1-1 downto 0 );
    q_13 : out std_logic_vector( 1-1 downto 0 );
    q_14 : out std_logic_vector( 1-1 downto 0 );
    q_15 : out std_logic_vector( 1-1 downto 0 );
    q_16 : out std_logic_vector( 1-1 downto 0 )
  );
end psb3_0_vector_delay_x5;
architecture structural of psb3_0_vector_delay_x5 is 
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay9_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay7_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay0_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay14_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay15_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay10_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay11_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay13_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay12_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal slice2_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal slice0_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 1-1 downto 0 );
begin
  q_1 <= delay0_q_net;
  q_2 <= delay1_q_net;
  q_3 <= delay2_q_net;
  q_4 <= delay3_q_net;
  q_5 <= delay4_q_net;
  q_6 <= delay5_q_net;
  q_7 <= delay6_q_net;
  q_8 <= delay7_q_net;
  q_9 <= delay8_q_net;
  q_10 <= delay9_q_net;
  q_11 <= delay10_q_net;
  q_12 <= delay11_q_net;
  q_13 <= delay12_q_net;
  q_14 <= delay13_q_net;
  q_15 <= delay14_q_net;
  q_16 <= delay15_q_net;
  slice0_y_net <= d_1;
  slice1_y_net <= d_2;
  slice2_y_net <= d_3;
  slice3_y_net <= d_4;
  slice4_y_net <= d_5;
  slice5_y_net <= d_6;
  slice6_y_net <= d_7;
  slice7_y_net <= d_8;
  slice8_y_net <= d_9;
  slice9_y_net <= d_10;
  slice10_y_net <= d_11;
  slice11_y_net <= d_12;
  slice12_y_net <= d_13;
  slice13_y_net <= d_14;
  slice14_y_net <= d_15;
  slice15_y_net <= d_16;
  clk_net <= clk_1;
  ce_net <= ce_1;
  delay0 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice0_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay0_q_net
  );
  delay1 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice2_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay3 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice3_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  delay4 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice4_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net
  );
  delay5 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice5_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  delay6 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice6_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay6_q_net
  );
  delay7 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice7_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay7_q_net
  );
  delay8 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice8_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay8_q_net
  );
  delay9 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice9_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay9_q_net
  );
  delay10 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice10_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay10_q_net
  );
  delay11 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice11_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay11_q_net
  );
  delay12 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice12_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay12_q_net
  );
  delay13 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice13_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay13_q_net
  );
  delay14 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice14_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay14_q_net
  );
  delay15 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice15_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay15_q_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Overflow Detector add_re_3/Vector Delay1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_delay1_x5 is
  port (
    d_1 : in std_logic_vector( 1-1 downto 0 );
    d_2 : in std_logic_vector( 1-1 downto 0 );
    d_3 : in std_logic_vector( 1-1 downto 0 );
    d_4 : in std_logic_vector( 1-1 downto 0 );
    d_5 : in std_logic_vector( 1-1 downto 0 );
    d_6 : in std_logic_vector( 1-1 downto 0 );
    d_7 : in std_logic_vector( 1-1 downto 0 );
    d_8 : in std_logic_vector( 1-1 downto 0 );
    d_9 : in std_logic_vector( 1-1 downto 0 );
    d_10 : in std_logic_vector( 1-1 downto 0 );
    d_11 : in std_logic_vector( 1-1 downto 0 );
    d_12 : in std_logic_vector( 1-1 downto 0 );
    d_13 : in std_logic_vector( 1-1 downto 0 );
    d_14 : in std_logic_vector( 1-1 downto 0 );
    d_15 : in std_logic_vector( 1-1 downto 0 );
    d_16 : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    q_1 : out std_logic_vector( 1-1 downto 0 );
    q_2 : out std_logic_vector( 1-1 downto 0 );
    q_3 : out std_logic_vector( 1-1 downto 0 );
    q_4 : out std_logic_vector( 1-1 downto 0 );
    q_5 : out std_logic_vector( 1-1 downto 0 );
    q_6 : out std_logic_vector( 1-1 downto 0 );
    q_7 : out std_logic_vector( 1-1 downto 0 );
    q_8 : out std_logic_vector( 1-1 downto 0 );
    q_9 : out std_logic_vector( 1-1 downto 0 );
    q_10 : out std_logic_vector( 1-1 downto 0 );
    q_11 : out std_logic_vector( 1-1 downto 0 );
    q_12 : out std_logic_vector( 1-1 downto 0 );
    q_13 : out std_logic_vector( 1-1 downto 0 );
    q_14 : out std_logic_vector( 1-1 downto 0 );
    q_15 : out std_logic_vector( 1-1 downto 0 );
    q_16 : out std_logic_vector( 1-1 downto 0 )
  );
end psb3_0_vector_delay1_x5;
architecture structural of psb3_0_vector_delay1_x5 is 
  signal slice6_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay15_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay14_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay13_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay11_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay0_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay7_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay9_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay10_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay12_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal slice15_y_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
begin
  q_1 <= delay0_q_net;
  q_2 <= delay1_q_net;
  q_3 <= delay2_q_net;
  q_4 <= delay3_q_net;
  q_5 <= delay4_q_net;
  q_6 <= delay5_q_net;
  q_7 <= delay6_q_net;
  q_8 <= delay7_q_net;
  q_9 <= delay8_q_net;
  q_10 <= delay9_q_net;
  q_11 <= delay10_q_net;
  q_12 <= delay11_q_net;
  q_13 <= delay12_q_net;
  q_14 <= delay13_q_net;
  q_15 <= delay14_q_net;
  q_16 <= delay15_q_net;
  slice0_y_net <= d_1;
  slice1_y_net <= d_2;
  slice2_y_net <= d_3;
  slice3_y_net <= d_4;
  slice4_y_net <= d_5;
  slice5_y_net <= d_6;
  slice6_y_net <= d_7;
  slice7_y_net <= d_8;
  slice8_y_net <= d_9;
  slice9_y_net <= d_10;
  slice10_y_net <= d_11;
  slice11_y_net <= d_12;
  slice12_y_net <= d_13;
  slice13_y_net <= d_14;
  slice14_y_net <= d_15;
  slice15_y_net <= d_16;
  clk_net <= clk_1;
  ce_net <= ce_1;
  delay0 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice0_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay0_q_net
  );
  delay1 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice2_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay3 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice3_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  delay4 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice4_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net
  );
  delay5 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice5_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  delay6 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice6_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay6_q_net
  );
  delay7 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice7_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay7_q_net
  );
  delay8 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice8_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay8_q_net
  );
  delay9 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice9_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay9_q_net
  );
  delay10 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice10_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay10_q_net
  );
  delay11 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice11_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay11_q_net
  );
  delay12 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice12_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay12_q_net
  );
  delay13 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice13_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay13_q_net
  );
  delay14 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice14_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay14_q_net
  );
  delay15 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice15_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay15_q_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Overflow Detector add_re_3/Vector Slice
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_slice_x5 is
  port (
    in_1 : in std_logic_vector( 16-1 downto 0 );
    in_2 : in std_logic_vector( 16-1 downto 0 );
    in_3 : in std_logic_vector( 16-1 downto 0 );
    in_4 : in std_logic_vector( 16-1 downto 0 );
    in_5 : in std_logic_vector( 16-1 downto 0 );
    in_6 : in std_logic_vector( 16-1 downto 0 );
    in_7 : in std_logic_vector( 16-1 downto 0 );
    in_8 : in std_logic_vector( 16-1 downto 0 );
    in_9 : in std_logic_vector( 16-1 downto 0 );
    in_10 : in std_logic_vector( 16-1 downto 0 );
    in_11 : in std_logic_vector( 16-1 downto 0 );
    in_12 : in std_logic_vector( 16-1 downto 0 );
    in_13 : in std_logic_vector( 16-1 downto 0 );
    in_14 : in std_logic_vector( 16-1 downto 0 );
    in_15 : in std_logic_vector( 16-1 downto 0 );
    in_16 : in std_logic_vector( 16-1 downto 0 );
    out_1 : out std_logic_vector( 1-1 downto 0 );
    out_2 : out std_logic_vector( 1-1 downto 0 );
    out_3 : out std_logic_vector( 1-1 downto 0 );
    out_4 : out std_logic_vector( 1-1 downto 0 );
    out_5 : out std_logic_vector( 1-1 downto 0 );
    out_6 : out std_logic_vector( 1-1 downto 0 );
    out_7 : out std_logic_vector( 1-1 downto 0 );
    out_8 : out std_logic_vector( 1-1 downto 0 );
    out_9 : out std_logic_vector( 1-1 downto 0 );
    out_10 : out std_logic_vector( 1-1 downto 0 );
    out_11 : out std_logic_vector( 1-1 downto 0 );
    out_12 : out std_logic_vector( 1-1 downto 0 );
    out_13 : out std_logic_vector( 1-1 downto 0 );
    out_14 : out std_logic_vector( 1-1 downto 0 );
    out_15 : out std_logic_vector( 1-1 downto 0 );
    out_16 : out std_logic_vector( 1-1 downto 0 )
  );
end psb3_0_vector_slice_x5;
architecture structural of psb3_0_vector_slice_x5 is 
  signal slice1_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 1-1 downto 0 );
  signal mult10_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult7_p_net : std_logic_vector( 16-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 1-1 downto 0 );
  signal mult14_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult2_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult9_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult8_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult11_p_net : std_logic_vector( 16-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 1-1 downto 0 );
  signal mult0_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult12_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult1_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult4_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult13_p_net : std_logic_vector( 16-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 1-1 downto 0 );
  signal mult5_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult6_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult3_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult15_p_net : std_logic_vector( 16-1 downto 0 );
begin
  out_1 <= slice0_y_net;
  out_2 <= slice1_y_net;
  out_3 <= slice2_y_net;
  out_4 <= slice3_y_net;
  out_5 <= slice4_y_net;
  out_6 <= slice5_y_net;
  out_7 <= slice6_y_net;
  out_8 <= slice7_y_net;
  out_9 <= slice8_y_net;
  out_10 <= slice9_y_net;
  out_11 <= slice10_y_net;
  out_12 <= slice11_y_net;
  out_13 <= slice12_y_net;
  out_14 <= slice13_y_net;
  out_15 <= slice14_y_net;
  out_16 <= slice15_y_net;
  mult0_p_net <= in_1;
  mult1_p_net <= in_2;
  mult2_p_net <= in_3;
  mult3_p_net <= in_4;
  mult4_p_net <= in_5;
  mult5_p_net <= in_6;
  mult6_p_net <= in_7;
  mult7_p_net <= in_8;
  mult8_p_net <= in_9;
  mult9_p_net <= in_10;
  mult10_p_net <= in_11;
  mult11_p_net <= in_12;
  mult12_p_net <= in_13;
  mult13_p_net <= in_14;
  mult14_p_net <= in_15;
  mult15_p_net <= in_16;
  slice0 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult0_p_net,
    y => slice0_y_net
  );
  slice1 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult1_p_net,
    y => slice1_y_net
  );
  slice2 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult2_p_net,
    y => slice2_y_net
  );
  slice3 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult3_p_net,
    y => slice3_y_net
  );
  slice4 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult4_p_net,
    y => slice4_y_net
  );
  slice5 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult5_p_net,
    y => slice5_y_net
  );
  slice6 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult6_p_net,
    y => slice6_y_net
  );
  slice7 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult7_p_net,
    y => slice7_y_net
  );
  slice8 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult8_p_net,
    y => slice8_y_net
  );
  slice9 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult9_p_net,
    y => slice9_y_net
  );
  slice10 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult10_p_net,
    y => slice10_y_net
  );
  slice11 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult11_p_net,
    y => slice11_y_net
  );
  slice12 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult12_p_net,
    y => slice12_y_net
  );
  slice13 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult13_p_net,
    y => slice13_y_net
  );
  slice14 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult14_p_net,
    y => slice14_y_net
  );
  slice15 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult15_p_net,
    y => slice15_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Overflow Detector add_re_3/Vector Slice1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_slice1_x5 is
  port (
    in_1 : in std_logic_vector( 16-1 downto 0 );
    in_2 : in std_logic_vector( 16-1 downto 0 );
    in_3 : in std_logic_vector( 16-1 downto 0 );
    in_4 : in std_logic_vector( 16-1 downto 0 );
    in_5 : in std_logic_vector( 16-1 downto 0 );
    in_6 : in std_logic_vector( 16-1 downto 0 );
    in_7 : in std_logic_vector( 16-1 downto 0 );
    in_8 : in std_logic_vector( 16-1 downto 0 );
    in_9 : in std_logic_vector( 16-1 downto 0 );
    in_10 : in std_logic_vector( 16-1 downto 0 );
    in_11 : in std_logic_vector( 16-1 downto 0 );
    in_12 : in std_logic_vector( 16-1 downto 0 );
    in_13 : in std_logic_vector( 16-1 downto 0 );
    in_14 : in std_logic_vector( 16-1 downto 0 );
    in_15 : in std_logic_vector( 16-1 downto 0 );
    in_16 : in std_logic_vector( 16-1 downto 0 );
    out_1 : out std_logic_vector( 1-1 downto 0 );
    out_2 : out std_logic_vector( 1-1 downto 0 );
    out_3 : out std_logic_vector( 1-1 downto 0 );
    out_4 : out std_logic_vector( 1-1 downto 0 );
    out_5 : out std_logic_vector( 1-1 downto 0 );
    out_6 : out std_logic_vector( 1-1 downto 0 );
    out_7 : out std_logic_vector( 1-1 downto 0 );
    out_8 : out std_logic_vector( 1-1 downto 0 );
    out_9 : out std_logic_vector( 1-1 downto 0 );
    out_10 : out std_logic_vector( 1-1 downto 0 );
    out_11 : out std_logic_vector( 1-1 downto 0 );
    out_12 : out std_logic_vector( 1-1 downto 0 );
    out_13 : out std_logic_vector( 1-1 downto 0 );
    out_14 : out std_logic_vector( 1-1 downto 0 );
    out_15 : out std_logic_vector( 1-1 downto 0 );
    out_16 : out std_logic_vector( 1-1 downto 0 )
  );
end psb3_0_vector_slice1_x5;
architecture structural of psb3_0_vector_slice1_x5 is 
  signal slice12_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
begin
  out_1 <= slice0_y_net;
  out_2 <= slice1_y_net;
  out_3 <= slice2_y_net;
  out_4 <= slice3_y_net;
  out_5 <= slice4_y_net;
  out_6 <= slice5_y_net;
  out_7 <= slice6_y_net;
  out_8 <= slice7_y_net;
  out_9 <= slice8_y_net;
  out_10 <= slice9_y_net;
  out_11 <= slice10_y_net;
  out_12 <= slice11_y_net;
  out_13 <= slice12_y_net;
  out_14 <= slice13_y_net;
  out_15 <= slice14_y_net;
  out_16 <= slice15_y_net;
  reinterpret0_output_port_net <= in_1;
  reinterpret1_output_port_net <= in_2;
  reinterpret2_output_port_net <= in_3;
  reinterpret3_output_port_net <= in_4;
  reinterpret4_output_port_net <= in_5;
  reinterpret5_output_port_net <= in_6;
  reinterpret6_output_port_net <= in_7;
  reinterpret7_output_port_net <= in_8;
  reinterpret8_output_port_net <= in_9;
  reinterpret9_output_port_net <= in_10;
  reinterpret10_output_port_net <= in_11;
  reinterpret11_output_port_net <= in_12;
  reinterpret12_output_port_net <= in_13;
  reinterpret13_output_port_net <= in_14;
  reinterpret14_output_port_net <= in_15;
  reinterpret15_output_port_net <= in_16;
  slice0 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret0_output_port_net,
    y => slice0_y_net
  );
  slice1 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret1_output_port_net,
    y => slice1_y_net
  );
  slice2 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret2_output_port_net,
    y => slice2_y_net
  );
  slice3 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret3_output_port_net,
    y => slice3_y_net
  );
  slice4 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret4_output_port_net,
    y => slice4_y_net
  );
  slice5 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret5_output_port_net,
    y => slice5_y_net
  );
  slice6 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret6_output_port_net,
    y => slice6_y_net
  );
  slice7 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret7_output_port_net,
    y => slice7_y_net
  );
  slice8 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret8_output_port_net,
    y => slice8_y_net
  );
  slice9 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret9_output_port_net,
    y => slice9_y_net
  );
  slice10 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret10_output_port_net,
    y => slice10_y_net
  );
  slice11 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret11_output_port_net,
    y => slice11_y_net
  );
  slice12 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret12_output_port_net,
    y => slice12_y_net
  );
  slice13 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret13_output_port_net,
    y => slice13_y_net
  );
  slice14 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret14_output_port_net,
    y => slice14_y_net
  );
  slice15 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret15_output_port_net,
    y => slice15_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Overflow Detector add_re_3/Vector Slice2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_slice2_x5 is
  port (
    in_1 : in std_logic_vector( 16-1 downto 0 );
    in_2 : in std_logic_vector( 16-1 downto 0 );
    in_3 : in std_logic_vector( 16-1 downto 0 );
    in_4 : in std_logic_vector( 16-1 downto 0 );
    in_5 : in std_logic_vector( 16-1 downto 0 );
    in_6 : in std_logic_vector( 16-1 downto 0 );
    in_7 : in std_logic_vector( 16-1 downto 0 );
    in_8 : in std_logic_vector( 16-1 downto 0 );
    in_9 : in std_logic_vector( 16-1 downto 0 );
    in_10 : in std_logic_vector( 16-1 downto 0 );
    in_11 : in std_logic_vector( 16-1 downto 0 );
    in_12 : in std_logic_vector( 16-1 downto 0 );
    in_13 : in std_logic_vector( 16-1 downto 0 );
    in_14 : in std_logic_vector( 16-1 downto 0 );
    in_15 : in std_logic_vector( 16-1 downto 0 );
    in_16 : in std_logic_vector( 16-1 downto 0 );
    out_1 : out std_logic_vector( 1-1 downto 0 );
    out_2 : out std_logic_vector( 1-1 downto 0 );
    out_3 : out std_logic_vector( 1-1 downto 0 );
    out_4 : out std_logic_vector( 1-1 downto 0 );
    out_5 : out std_logic_vector( 1-1 downto 0 );
    out_6 : out std_logic_vector( 1-1 downto 0 );
    out_7 : out std_logic_vector( 1-1 downto 0 );
    out_8 : out std_logic_vector( 1-1 downto 0 );
    out_9 : out std_logic_vector( 1-1 downto 0 );
    out_10 : out std_logic_vector( 1-1 downto 0 );
    out_11 : out std_logic_vector( 1-1 downto 0 );
    out_12 : out std_logic_vector( 1-1 downto 0 );
    out_13 : out std_logic_vector( 1-1 downto 0 );
    out_14 : out std_logic_vector( 1-1 downto 0 );
    out_15 : out std_logic_vector( 1-1 downto 0 );
    out_16 : out std_logic_vector( 1-1 downto 0 )
  );
end psb3_0_vector_slice2_x5;
architecture structural of psb3_0_vector_slice2_x5 is 
  signal addsub0_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub3_s_net : std_logic_vector( 16-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 1-1 downto 0 );
  signal addsub7_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub11_s_net : std_logic_vector( 16-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 1-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 16-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 1-1 downto 0 );
  signal addsub8_s_net : std_logic_vector( 16-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 1-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub9_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub12_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub14_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub6_s_net : std_logic_vector( 16-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 1-1 downto 0 );
  signal addsub13_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub5_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub10_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub15_s_net : std_logic_vector( 16-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 1-1 downto 0 );
begin
  out_1 <= slice0_y_net;
  out_2 <= slice1_y_net;
  out_3 <= slice2_y_net;
  out_4 <= slice3_y_net;
  out_5 <= slice4_y_net;
  out_6 <= slice5_y_net;
  out_7 <= slice6_y_net;
  out_8 <= slice7_y_net;
  out_9 <= slice8_y_net;
  out_10 <= slice9_y_net;
  out_11 <= slice10_y_net;
  out_12 <= slice11_y_net;
  out_13 <= slice12_y_net;
  out_14 <= slice13_y_net;
  out_15 <= slice14_y_net;
  out_16 <= slice15_y_net;
  addsub0_s_net <= in_1;
  addsub1_s_net <= in_2;
  addsub2_s_net <= in_3;
  addsub3_s_net <= in_4;
  addsub4_s_net <= in_5;
  addsub5_s_net <= in_6;
  addsub6_s_net <= in_7;
  addsub7_s_net <= in_8;
  addsub8_s_net <= in_9;
  addsub9_s_net <= in_10;
  addsub10_s_net <= in_11;
  addsub11_s_net <= in_12;
  addsub12_s_net <= in_13;
  addsub13_s_net <= in_14;
  addsub14_s_net <= in_15;
  addsub15_s_net <= in_16;
  slice0 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub0_s_net,
    y => slice0_y_net
  );
  slice1 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub1_s_net,
    y => slice1_y_net
  );
  slice2 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub2_s_net,
    y => slice2_y_net
  );
  slice3 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub3_s_net,
    y => slice3_y_net
  );
  slice4 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub4_s_net,
    y => slice4_y_net
  );
  slice5 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub5_s_net,
    y => slice5_y_net
  );
  slice6 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub6_s_net,
    y => slice6_y_net
  );
  slice7 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub7_s_net,
    y => slice7_y_net
  );
  slice8 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub8_s_net,
    y => slice8_y_net
  );
  slice9 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub9_s_net,
    y => slice9_y_net
  );
  slice10 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub10_s_net,
    y => slice10_y_net
  );
  slice11 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub11_s_net,
    y => slice11_y_net
  );
  slice12 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub12_s_net,
    y => slice12_y_net
  );
  slice13 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub13_s_net,
    y => slice13_y_net
  );
  slice14 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub14_s_net,
    y => slice14_y_net
  );
  slice15 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub15_s_net,
    y => slice15_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Overflow Detector add_re_3/Vector to Scalar
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_to_scalar_x5 is
  port (
    i_1 : in std_logic_vector( 1-1 downto 0 );
    i_2 : in std_logic_vector( 1-1 downto 0 );
    i_3 : in std_logic_vector( 1-1 downto 0 );
    i_4 : in std_logic_vector( 1-1 downto 0 );
    i_5 : in std_logic_vector( 1-1 downto 0 );
    i_6 : in std_logic_vector( 1-1 downto 0 );
    i_7 : in std_logic_vector( 1-1 downto 0 );
    i_8 : in std_logic_vector( 1-1 downto 0 );
    i_9 : in std_logic_vector( 1-1 downto 0 );
    i_10 : in std_logic_vector( 1-1 downto 0 );
    i_11 : in std_logic_vector( 1-1 downto 0 );
    i_12 : in std_logic_vector( 1-1 downto 0 );
    i_13 : in std_logic_vector( 1-1 downto 0 );
    i_14 : in std_logic_vector( 1-1 downto 0 );
    i_15 : in std_logic_vector( 1-1 downto 0 );
    i_16 : in std_logic_vector( 1-1 downto 0 );
    o : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_vector_to_scalar_x5;
architecture structural of psb3_0_vector_to_scalar_x5 is 
  signal delay15_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay10_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay7_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay14_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay11_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay12_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal concat1_y_net : std_logic_vector( 16-1 downto 0 );
  signal delay0_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay9_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay13_q_net : std_logic_vector( 1-1 downto 0 );
begin
  o <= concat1_y_net;
  delay0_q_net <= i_1;
  delay1_q_net <= i_2;
  delay2_q_net <= i_3;
  delay3_q_net <= i_4;
  delay4_q_net <= i_5;
  delay5_q_net <= i_6;
  delay6_q_net <= i_7;
  delay7_q_net <= i_8;
  delay8_q_net <= i_9;
  delay9_q_net <= i_10;
  delay10_q_net <= i_11;
  delay11_q_net <= i_12;
  delay12_q_net <= i_13;
  delay13_q_net <= i_14;
  delay14_q_net <= i_15;
  delay15_q_net <= i_16;
  concat1 : entity xil_defaultlib.sysgen_concat_d977c66e35 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => delay15_q_net,
    in1 => delay14_q_net,
    in2 => delay13_q_net,
    in3 => delay12_q_net,
    in4 => delay11_q_net,
    in5 => delay10_q_net,
    in6 => delay9_q_net,
    in7 => delay8_q_net,
    in8 => delay7_q_net,
    in9 => delay6_q_net,
    in10 => delay5_q_net,
    in11 => delay4_q_net,
    in12 => delay3_q_net,
    in13 => delay2_q_net,
    in14 => delay1_q_net,
    in15 => delay0_q_net,
    y => concat1_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Overflow Detector add_re_3/Vector to Scalar1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_to_scalar1_x5 is
  port (
    i_1 : in std_logic_vector( 1-1 downto 0 );
    i_2 : in std_logic_vector( 1-1 downto 0 );
    i_3 : in std_logic_vector( 1-1 downto 0 );
    i_4 : in std_logic_vector( 1-1 downto 0 );
    i_5 : in std_logic_vector( 1-1 downto 0 );
    i_6 : in std_logic_vector( 1-1 downto 0 );
    i_7 : in std_logic_vector( 1-1 downto 0 );
    i_8 : in std_logic_vector( 1-1 downto 0 );
    i_9 : in std_logic_vector( 1-1 downto 0 );
    i_10 : in std_logic_vector( 1-1 downto 0 );
    i_11 : in std_logic_vector( 1-1 downto 0 );
    i_12 : in std_logic_vector( 1-1 downto 0 );
    i_13 : in std_logic_vector( 1-1 downto 0 );
    i_14 : in std_logic_vector( 1-1 downto 0 );
    i_15 : in std_logic_vector( 1-1 downto 0 );
    i_16 : in std_logic_vector( 1-1 downto 0 );
    o : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_vector_to_scalar1_x5;
architecture structural of psb3_0_vector_to_scalar1_x5 is 
  signal delay12_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay14_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay10_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay0_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay11_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay15_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay9_q_net : std_logic_vector( 1-1 downto 0 );
  signal concat1_y_net : std_logic_vector( 16-1 downto 0 );
  signal delay13_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay7_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 1-1 downto 0 );
begin
  o <= concat1_y_net;
  delay0_q_net <= i_1;
  delay1_q_net <= i_2;
  delay2_q_net <= i_3;
  delay3_q_net <= i_4;
  delay4_q_net <= i_5;
  delay5_q_net <= i_6;
  delay6_q_net <= i_7;
  delay7_q_net <= i_8;
  delay8_q_net <= i_9;
  delay9_q_net <= i_10;
  delay10_q_net <= i_11;
  delay11_q_net <= i_12;
  delay12_q_net <= i_13;
  delay13_q_net <= i_14;
  delay14_q_net <= i_15;
  delay15_q_net <= i_16;
  concat1 : entity xil_defaultlib.sysgen_concat_d977c66e35 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => delay15_q_net,
    in1 => delay14_q_net,
    in2 => delay13_q_net,
    in3 => delay12_q_net,
    in4 => delay11_q_net,
    in5 => delay10_q_net,
    in6 => delay9_q_net,
    in7 => delay8_q_net,
    in8 => delay7_q_net,
    in9 => delay6_q_net,
    in10 => delay5_q_net,
    in11 => delay4_q_net,
    in12 => delay3_q_net,
    in13 => delay2_q_net,
    in14 => delay1_q_net,
    in15 => delay0_q_net,
    y => concat1_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Overflow Detector add_re_3/Vector to Scalar2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_to_scalar2_x5 is
  port (
    i_1 : in std_logic_vector( 1-1 downto 0 );
    i_2 : in std_logic_vector( 1-1 downto 0 );
    i_3 : in std_logic_vector( 1-1 downto 0 );
    i_4 : in std_logic_vector( 1-1 downto 0 );
    i_5 : in std_logic_vector( 1-1 downto 0 );
    i_6 : in std_logic_vector( 1-1 downto 0 );
    i_7 : in std_logic_vector( 1-1 downto 0 );
    i_8 : in std_logic_vector( 1-1 downto 0 );
    i_9 : in std_logic_vector( 1-1 downto 0 );
    i_10 : in std_logic_vector( 1-1 downto 0 );
    i_11 : in std_logic_vector( 1-1 downto 0 );
    i_12 : in std_logic_vector( 1-1 downto 0 );
    i_13 : in std_logic_vector( 1-1 downto 0 );
    i_14 : in std_logic_vector( 1-1 downto 0 );
    i_15 : in std_logic_vector( 1-1 downto 0 );
    i_16 : in std_logic_vector( 1-1 downto 0 );
    o : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_vector_to_scalar2_x5;
architecture structural of psb3_0_vector_to_scalar2_x5 is 
  signal slice5_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 1-1 downto 0 );
  signal concat1_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 1-1 downto 0 );
begin
  o <= concat1_y_net;
  slice0_y_net <= i_1;
  slice1_y_net <= i_2;
  slice2_y_net <= i_3;
  slice3_y_net <= i_4;
  slice4_y_net <= i_5;
  slice5_y_net <= i_6;
  slice6_y_net <= i_7;
  slice7_y_net <= i_8;
  slice8_y_net <= i_9;
  slice9_y_net <= i_10;
  slice10_y_net <= i_11;
  slice11_y_net <= i_12;
  slice12_y_net <= i_13;
  slice13_y_net <= i_14;
  slice14_y_net <= i_15;
  slice15_y_net <= i_16;
  concat1 : entity xil_defaultlib.sysgen_concat_d977c66e35 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => slice15_y_net,
    in1 => slice14_y_net,
    in2 => slice13_y_net,
    in3 => slice12_y_net,
    in4 => slice11_y_net,
    in5 => slice10_y_net,
    in6 => slice9_y_net,
    in7 => slice8_y_net,
    in8 => slice7_y_net,
    in9 => slice6_y_net,
    in10 => slice5_y_net,
    in11 => slice4_y_net,
    in12 => slice3_y_net,
    in13 => slice2_y_net,
    in14 => slice1_y_net,
    in15 => slice0_y_net,
    y => concat1_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Overflow Detector add_re_3
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_overflow_detector_add_re_3 is
  port (
    rst : in std_logic_vector( 1-1 downto 0 );
    a_1 : in std_logic_vector( 16-1 downto 0 );
    b_1 : in std_logic_vector( 16-1 downto 0 );
    s_1 : in std_logic_vector( 16-1 downto 0 );
    a_2 : in std_logic_vector( 16-1 downto 0 );
    a_3 : in std_logic_vector( 16-1 downto 0 );
    a_4 : in std_logic_vector( 16-1 downto 0 );
    a_5 : in std_logic_vector( 16-1 downto 0 );
    a_6 : in std_logic_vector( 16-1 downto 0 );
    a_7 : in std_logic_vector( 16-1 downto 0 );
    a_8 : in std_logic_vector( 16-1 downto 0 );
    a_9 : in std_logic_vector( 16-1 downto 0 );
    a_10 : in std_logic_vector( 16-1 downto 0 );
    a_11 : in std_logic_vector( 16-1 downto 0 );
    a_12 : in std_logic_vector( 16-1 downto 0 );
    a_13 : in std_logic_vector( 16-1 downto 0 );
    a_14 : in std_logic_vector( 16-1 downto 0 );
    a_15 : in std_logic_vector( 16-1 downto 0 );
    a_16 : in std_logic_vector( 16-1 downto 0 );
    b_2 : in std_logic_vector( 16-1 downto 0 );
    b_3 : in std_logic_vector( 16-1 downto 0 );
    b_4 : in std_logic_vector( 16-1 downto 0 );
    b_5 : in std_logic_vector( 16-1 downto 0 );
    b_6 : in std_logic_vector( 16-1 downto 0 );
    b_7 : in std_logic_vector( 16-1 downto 0 );
    b_8 : in std_logic_vector( 16-1 downto 0 );
    b_9 : in std_logic_vector( 16-1 downto 0 );
    b_10 : in std_logic_vector( 16-1 downto 0 );
    b_11 : in std_logic_vector( 16-1 downto 0 );
    b_12 : in std_logic_vector( 16-1 downto 0 );
    b_13 : in std_logic_vector( 16-1 downto 0 );
    b_14 : in std_logic_vector( 16-1 downto 0 );
    b_15 : in std_logic_vector( 16-1 downto 0 );
    b_16 : in std_logic_vector( 16-1 downto 0 );
    s_2 : in std_logic_vector( 16-1 downto 0 );
    s_3 : in std_logic_vector( 16-1 downto 0 );
    s_4 : in std_logic_vector( 16-1 downto 0 );
    s_5 : in std_logic_vector( 16-1 downto 0 );
    s_6 : in std_logic_vector( 16-1 downto 0 );
    s_7 : in std_logic_vector( 16-1 downto 0 );
    s_8 : in std_logic_vector( 16-1 downto 0 );
    s_9 : in std_logic_vector( 16-1 downto 0 );
    s_10 : in std_logic_vector( 16-1 downto 0 );
    s_11 : in std_logic_vector( 16-1 downto 0 );
    s_12 : in std_logic_vector( 16-1 downto 0 );
    s_13 : in std_logic_vector( 16-1 downto 0 );
    s_14 : in std_logic_vector( 16-1 downto 0 );
    s_15 : in std_logic_vector( 16-1 downto 0 );
    s_16 : in std_logic_vector( 16-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    ov : out std_logic_vector( 1-1 downto 0 )
  );
end psb3_0_overflow_detector_add_re_3;
architecture structural of psb3_0_overflow_detector_add_re_3 is 
  signal register_q_net : std_logic_vector( 1-1 downto 0 );
  signal gin_tl_reset_net : std_logic_vector( 1-1 downto 0 );
  signal mult0_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult15_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mult8_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mult7_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult11_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult9_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult12_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult13_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub0_s_net : std_logic_vector( 16-1 downto 0 );
  signal mult4_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult1_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mult2_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult5_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mult6_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult14_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mult3_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult10_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub8_s_net : std_logic_vector( 16-1 downto 0 );
  signal delay2_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub7_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub14_s_net : std_logic_vector( 16-1 downto 0 );
  signal delay3_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay8_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal addsub11_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub10_s_net : std_logic_vector( 16-1 downto 0 );
  signal delay10_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice0_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 16-1 downto 0 );
  signal delay14_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice2_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal slice3_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal slice7_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 16-1 downto 0 );
  signal delay1_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay15_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice6_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal slice9_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal delay0_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal addsub12_s_net : std_logic_vector( 16-1 downto 0 );
  signal delay9_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay11_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay12_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay13_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice11_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal slice12_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal addsub5_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub6_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub9_s_net : std_logic_vector( 16-1 downto 0 );
  signal delay7_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal delay4_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal addsub13_s_net : std_logic_vector( 16-1 downto 0 );
  signal delay6_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice1_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal slice8_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal addsub3_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub15_s_net : std_logic_vector( 16-1 downto 0 );
  signal slice4_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal slice10_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal delay5_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal slice5_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice3_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 1-1 downto 0 );
  signal concat1_y_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal slice1_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice0_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal constant17_op_net : std_logic_vector( 1-1 downto 0 );
  signal slice9_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice4_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice7_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice2_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay12_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay13_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay15_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice8_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice13_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice14_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice12_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice15_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay7_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice15_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal slice10_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay11_q_net : std_logic_vector( 1-1 downto 0 );
  signal concat1_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice6_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay14_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay9_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice5_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice14_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal delay0_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice11_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice13_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal delay10_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 1-1 downto 0 );
  signal concat1_y_net_x1 : std_logic_vector( 16-1 downto 0 );
  signal expression_dout_net : std_logic_vector( 1-1 downto 0 );
  signal convert_dout_net : std_logic_vector( 1-1 downto 0 );
begin
  ov <= register_q_net;
  gin_tl_reset_net <= rst;
  mult0_p_net <= a_1;
  reinterpret0_output_port_net <= b_1;
  addsub0_s_net <= s_1;
  mult1_p_net <= a_2;
  mult2_p_net <= a_3;
  mult3_p_net <= a_4;
  mult4_p_net <= a_5;
  mult5_p_net <= a_6;
  mult6_p_net <= a_7;
  mult7_p_net <= a_8;
  mult8_p_net <= a_9;
  mult9_p_net <= a_10;
  mult10_p_net <= a_11;
  mult11_p_net <= a_12;
  mult12_p_net <= a_13;
  mult13_p_net <= a_14;
  mult14_p_net <= a_15;
  mult15_p_net <= a_16;
  reinterpret1_output_port_net <= b_2;
  reinterpret2_output_port_net <= b_3;
  reinterpret3_output_port_net <= b_4;
  reinterpret4_output_port_net <= b_5;
  reinterpret5_output_port_net <= b_6;
  reinterpret6_output_port_net <= b_7;
  reinterpret7_output_port_net <= b_8;
  reinterpret8_output_port_net <= b_9;
  reinterpret9_output_port_net <= b_10;
  reinterpret10_output_port_net <= b_11;
  reinterpret11_output_port_net <= b_12;
  reinterpret12_output_port_net <= b_13;
  reinterpret13_output_port_net <= b_14;
  reinterpret14_output_port_net <= b_15;
  reinterpret15_output_port_net <= b_16;
  addsub1_s_net <= s_2;
  addsub2_s_net <= s_3;
  addsub3_s_net <= s_4;
  addsub4_s_net <= s_5;
  addsub5_s_net <= s_6;
  addsub6_s_net <= s_7;
  addsub7_s_net <= s_8;
  addsub8_s_net <= s_9;
  addsub9_s_net <= s_10;
  addsub10_s_net <= s_11;
  addsub11_s_net <= s_12;
  addsub12_s_net <= s_13;
  addsub13_s_net <= s_14;
  addsub14_s_net <= s_15;
  addsub15_s_net <= s_16;
  clk_net <= clk_1;
  ce_net <= ce_1;
  vector_delay : entity xil_defaultlib.psb3_0_vector_delay_x5 
  port map (
    d_1 => slice0_y_net_x1,
    d_2 => slice1_y_net_x1,
    d_3 => slice2_y_net_x1,
    d_4 => slice3_y_net_x1,
    d_5 => slice4_y_net_x1,
    d_6 => slice5_y_net_x1,
    d_7 => slice6_y_net_x1,
    d_8 => slice7_y_net_x1,
    d_9 => slice8_y_net_x1,
    d_10 => slice9_y_net_x1,
    d_11 => slice10_y_net_x1,
    d_12 => slice11_y_net_x1,
    d_13 => slice12_y_net_x1,
    d_14 => slice13_y_net_x1,
    d_15 => slice14_y_net_x1,
    d_16 => slice15_y_net_x1,
    clk_1 => clk_net,
    ce_1 => ce_net,
    q_1 => delay0_q_net_x0,
    q_2 => delay1_q_net_x0,
    q_3 => delay2_q_net_x0,
    q_4 => delay3_q_net_x0,
    q_5 => delay4_q_net_x0,
    q_6 => delay5_q_net_x0,
    q_7 => delay6_q_net_x0,
    q_8 => delay7_q_net_x0,
    q_9 => delay8_q_net_x0,
    q_10 => delay9_q_net_x0,
    q_11 => delay10_q_net_x0,
    q_12 => delay11_q_net_x0,
    q_13 => delay12_q_net_x0,
    q_14 => delay13_q_net_x0,
    q_15 => delay14_q_net_x0,
    q_16 => delay15_q_net_x0
  );
  vector_delay1 : entity xil_defaultlib.psb3_0_vector_delay1_x5 
  port map (
    d_1 => slice0_y_net_x0,
    d_2 => slice1_y_net_x0,
    d_3 => slice2_y_net_x0,
    d_4 => slice3_y_net_x0,
    d_5 => slice4_y_net_x0,
    d_6 => slice5_y_net_x0,
    d_7 => slice6_y_net_x0,
    d_8 => slice7_y_net_x0,
    d_9 => slice8_y_net_x0,
    d_10 => slice9_y_net_x0,
    d_11 => slice10_y_net_x0,
    d_12 => slice11_y_net_x0,
    d_13 => slice12_y_net_x0,
    d_14 => slice13_y_net_x0,
    d_15 => slice14_y_net_x0,
    d_16 => slice15_y_net_x0,
    clk_1 => clk_net,
    ce_1 => ce_net,
    q_1 => delay0_q_net,
    q_2 => delay1_q_net,
    q_3 => delay2_q_net,
    q_4 => delay3_q_net,
    q_5 => delay4_q_net,
    q_6 => delay5_q_net,
    q_7 => delay6_q_net,
    q_8 => delay7_q_net,
    q_9 => delay8_q_net,
    q_10 => delay9_q_net,
    q_11 => delay10_q_net,
    q_12 => delay11_q_net,
    q_13 => delay12_q_net,
    q_14 => delay13_q_net,
    q_15 => delay14_q_net,
    q_16 => delay15_q_net
  );
  vector_slice : entity xil_defaultlib.psb3_0_vector_slice_x5 
  port map (
    in_1 => mult0_p_net,
    in_2 => mult1_p_net,
    in_3 => mult2_p_net,
    in_4 => mult3_p_net,
    in_5 => mult4_p_net,
    in_6 => mult5_p_net,
    in_7 => mult6_p_net,
    in_8 => mult7_p_net,
    in_9 => mult8_p_net,
    in_10 => mult9_p_net,
    in_11 => mult10_p_net,
    in_12 => mult11_p_net,
    in_13 => mult12_p_net,
    in_14 => mult13_p_net,
    in_15 => mult14_p_net,
    in_16 => mult15_p_net,
    out_1 => slice0_y_net_x1,
    out_2 => slice1_y_net_x1,
    out_3 => slice2_y_net_x1,
    out_4 => slice3_y_net_x1,
    out_5 => slice4_y_net_x1,
    out_6 => slice5_y_net_x1,
    out_7 => slice6_y_net_x1,
    out_8 => slice7_y_net_x1,
    out_9 => slice8_y_net_x1,
    out_10 => slice9_y_net_x1,
    out_11 => slice10_y_net_x1,
    out_12 => slice11_y_net_x1,
    out_13 => slice12_y_net_x1,
    out_14 => slice13_y_net_x1,
    out_15 => slice14_y_net_x1,
    out_16 => slice15_y_net_x1
  );
  vector_slice1 : entity xil_defaultlib.psb3_0_vector_slice1_x5 
  port map (
    in_1 => reinterpret0_output_port_net,
    in_2 => reinterpret1_output_port_net,
    in_3 => reinterpret2_output_port_net,
    in_4 => reinterpret3_output_port_net,
    in_5 => reinterpret4_output_port_net,
    in_6 => reinterpret5_output_port_net,
    in_7 => reinterpret6_output_port_net,
    in_8 => reinterpret7_output_port_net,
    in_9 => reinterpret8_output_port_net,
    in_10 => reinterpret9_output_port_net,
    in_11 => reinterpret10_output_port_net,
    in_12 => reinterpret11_output_port_net,
    in_13 => reinterpret12_output_port_net,
    in_14 => reinterpret13_output_port_net,
    in_15 => reinterpret14_output_port_net,
    in_16 => reinterpret15_output_port_net,
    out_1 => slice0_y_net_x0,
    out_2 => slice1_y_net_x0,
    out_3 => slice2_y_net_x0,
    out_4 => slice3_y_net_x0,
    out_5 => slice4_y_net_x0,
    out_6 => slice5_y_net_x0,
    out_7 => slice6_y_net_x0,
    out_8 => slice7_y_net_x0,
    out_9 => slice8_y_net_x0,
    out_10 => slice9_y_net_x0,
    out_11 => slice10_y_net_x0,
    out_12 => slice11_y_net_x0,
    out_13 => slice12_y_net_x0,
    out_14 => slice13_y_net_x0,
    out_15 => slice14_y_net_x0,
    out_16 => slice15_y_net_x0
  );
  vector_slice2 : entity xil_defaultlib.psb3_0_vector_slice2_x5 
  port map (
    in_1 => addsub0_s_net,
    in_2 => addsub1_s_net,
    in_3 => addsub2_s_net,
    in_4 => addsub3_s_net,
    in_5 => addsub4_s_net,
    in_6 => addsub5_s_net,
    in_7 => addsub6_s_net,
    in_8 => addsub7_s_net,
    in_9 => addsub8_s_net,
    in_10 => addsub9_s_net,
    in_11 => addsub10_s_net,
    in_12 => addsub11_s_net,
    in_13 => addsub12_s_net,
    in_14 => addsub13_s_net,
    in_15 => addsub14_s_net,
    in_16 => addsub15_s_net,
    out_1 => slice0_y_net,
    out_2 => slice1_y_net,
    out_3 => slice2_y_net,
    out_4 => slice3_y_net,
    out_5 => slice4_y_net,
    out_6 => slice5_y_net,
    out_7 => slice6_y_net,
    out_8 => slice7_y_net,
    out_9 => slice8_y_net,
    out_10 => slice9_y_net,
    out_11 => slice10_y_net,
    out_12 => slice11_y_net,
    out_13 => slice12_y_net,
    out_14 => slice13_y_net,
    out_15 => slice14_y_net,
    out_16 => slice15_y_net
  );
  vector_to_scalar : entity xil_defaultlib.psb3_0_vector_to_scalar_x5 
  port map (
    i_1 => delay0_q_net_x0,
    i_2 => delay1_q_net_x0,
    i_3 => delay2_q_net_x0,
    i_4 => delay3_q_net_x0,
    i_5 => delay4_q_net_x0,
    i_6 => delay5_q_net_x0,
    i_7 => delay6_q_net_x0,
    i_8 => delay7_q_net_x0,
    i_9 => delay8_q_net_x0,
    i_10 => delay9_q_net_x0,
    i_11 => delay10_q_net_x0,
    i_12 => delay11_q_net_x0,
    i_13 => delay12_q_net_x0,
    i_14 => delay13_q_net_x0,
    i_15 => delay14_q_net_x0,
    i_16 => delay15_q_net_x0,
    o => concat1_y_net_x1
  );
  vector_to_scalar1 : entity xil_defaultlib.psb3_0_vector_to_scalar1_x5 
  port map (
    i_1 => delay0_q_net,
    i_2 => delay1_q_net,
    i_3 => delay2_q_net,
    i_4 => delay3_q_net,
    i_5 => delay4_q_net,
    i_6 => delay5_q_net,
    i_7 => delay6_q_net,
    i_8 => delay7_q_net,
    i_9 => delay8_q_net,
    i_10 => delay9_q_net,
    i_11 => delay10_q_net,
    i_12 => delay11_q_net,
    i_13 => delay12_q_net,
    i_14 => delay13_q_net,
    i_15 => delay14_q_net,
    i_16 => delay15_q_net,
    o => concat1_y_net_x0
  );
  vector_to_scalar2 : entity xil_defaultlib.psb3_0_vector_to_scalar2_x5 
  port map (
    i_1 => slice0_y_net,
    i_2 => slice1_y_net,
    i_3 => slice2_y_net,
    i_4 => slice3_y_net,
    i_5 => slice4_y_net,
    i_6 => slice5_y_net,
    i_7 => slice6_y_net,
    i_8 => slice7_y_net,
    i_9 => slice8_y_net,
    i_10 => slice9_y_net,
    i_11 => slice10_y_net,
    i_12 => slice11_y_net,
    i_13 => slice12_y_net,
    i_14 => slice13_y_net,
    i_15 => slice14_y_net,
    i_16 => slice15_y_net,
    o => concat1_y_net
  );
  constant17 : entity xil_defaultlib.sysgen_constant_71e89d757c 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant17_op_net
  );
  convert : entity xil_defaultlib.psb3_0_xlconvert 
  generic map (
    bool_conversion => 1,
    din_arith => 1,
    din_bin_pt => 0,
    din_width => 1,
    dout_arith => 1,
    dout_bin_pt => 0,
    dout_width => 1,
    latency => 1,
    overflow => xlWrap,
    quantization => xlTruncate
  )
  port map (
    clr => '0',
    en => "1",
    din => expression_dout_net,
    clk => clk_net,
    ce => ce_net,
    dout => convert_dout_net
  );
  expression : entity xil_defaultlib.sysgen_expr_7c83532765 
  port map (
    clr => '0',
    a => concat1_y_net_x1,
    b => concat1_y_net_x0,
    s => concat1_y_net,
    clk => clk_net,
    ce => ce_net,
    dout => expression_dout_net
  );
  register_x0 : entity xil_defaultlib.psb3_0_xlregister 
  generic map (
    d_width => 1,
    init_value => b"0"
  )
  port map (
    d => constant17_op_net,
    rst => gin_tl_reset_net,
    en => convert_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => register_q_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Overflow Detector add_re_4/Vector Delay
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_delay_x6 is
  port (
    d_1 : in std_logic_vector( 1-1 downto 0 );
    d_2 : in std_logic_vector( 1-1 downto 0 );
    d_3 : in std_logic_vector( 1-1 downto 0 );
    d_4 : in std_logic_vector( 1-1 downto 0 );
    d_5 : in std_logic_vector( 1-1 downto 0 );
    d_6 : in std_logic_vector( 1-1 downto 0 );
    d_7 : in std_logic_vector( 1-1 downto 0 );
    d_8 : in std_logic_vector( 1-1 downto 0 );
    d_9 : in std_logic_vector( 1-1 downto 0 );
    d_10 : in std_logic_vector( 1-1 downto 0 );
    d_11 : in std_logic_vector( 1-1 downto 0 );
    d_12 : in std_logic_vector( 1-1 downto 0 );
    d_13 : in std_logic_vector( 1-1 downto 0 );
    d_14 : in std_logic_vector( 1-1 downto 0 );
    d_15 : in std_logic_vector( 1-1 downto 0 );
    d_16 : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    q_1 : out std_logic_vector( 1-1 downto 0 );
    q_2 : out std_logic_vector( 1-1 downto 0 );
    q_3 : out std_logic_vector( 1-1 downto 0 );
    q_4 : out std_logic_vector( 1-1 downto 0 );
    q_5 : out std_logic_vector( 1-1 downto 0 );
    q_6 : out std_logic_vector( 1-1 downto 0 );
    q_7 : out std_logic_vector( 1-1 downto 0 );
    q_8 : out std_logic_vector( 1-1 downto 0 );
    q_9 : out std_logic_vector( 1-1 downto 0 );
    q_10 : out std_logic_vector( 1-1 downto 0 );
    q_11 : out std_logic_vector( 1-1 downto 0 );
    q_12 : out std_logic_vector( 1-1 downto 0 );
    q_13 : out std_logic_vector( 1-1 downto 0 );
    q_14 : out std_logic_vector( 1-1 downto 0 );
    q_15 : out std_logic_vector( 1-1 downto 0 );
    q_16 : out std_logic_vector( 1-1 downto 0 )
  );
end psb3_0_vector_delay_x6;
architecture structural of psb3_0_vector_delay_x6 is 
  signal delay3_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay13_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay11_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay15_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay14_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay10_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay7_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay12_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay0_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay9_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal slice10_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal slice12_y_net : std_logic_vector( 1-1 downto 0 );
begin
  q_1 <= delay0_q_net;
  q_2 <= delay1_q_net;
  q_3 <= delay2_q_net;
  q_4 <= delay3_q_net;
  q_5 <= delay4_q_net;
  q_6 <= delay5_q_net;
  q_7 <= delay6_q_net;
  q_8 <= delay7_q_net;
  q_9 <= delay8_q_net;
  q_10 <= delay9_q_net;
  q_11 <= delay10_q_net;
  q_12 <= delay11_q_net;
  q_13 <= delay12_q_net;
  q_14 <= delay13_q_net;
  q_15 <= delay14_q_net;
  q_16 <= delay15_q_net;
  slice0_y_net <= d_1;
  slice1_y_net <= d_2;
  slice2_y_net <= d_3;
  slice3_y_net <= d_4;
  slice4_y_net <= d_5;
  slice5_y_net <= d_6;
  slice6_y_net <= d_7;
  slice7_y_net <= d_8;
  slice8_y_net <= d_9;
  slice9_y_net <= d_10;
  slice10_y_net <= d_11;
  slice11_y_net <= d_12;
  slice12_y_net <= d_13;
  slice13_y_net <= d_14;
  slice14_y_net <= d_15;
  slice15_y_net <= d_16;
  clk_net <= clk_1;
  ce_net <= ce_1;
  delay0 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice0_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay0_q_net
  );
  delay1 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice2_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay3 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice3_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  delay4 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice4_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net
  );
  delay5 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice5_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  delay6 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice6_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay6_q_net
  );
  delay7 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice7_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay7_q_net
  );
  delay8 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice8_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay8_q_net
  );
  delay9 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice9_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay9_q_net
  );
  delay10 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice10_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay10_q_net
  );
  delay11 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice11_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay11_q_net
  );
  delay12 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice12_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay12_q_net
  );
  delay13 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice13_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay13_q_net
  );
  delay14 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice14_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay14_q_net
  );
  delay15 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice15_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay15_q_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Overflow Detector add_re_4/Vector Delay1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_delay1_x6 is
  port (
    d_1 : in std_logic_vector( 1-1 downto 0 );
    d_2 : in std_logic_vector( 1-1 downto 0 );
    d_3 : in std_logic_vector( 1-1 downto 0 );
    d_4 : in std_logic_vector( 1-1 downto 0 );
    d_5 : in std_logic_vector( 1-1 downto 0 );
    d_6 : in std_logic_vector( 1-1 downto 0 );
    d_7 : in std_logic_vector( 1-1 downto 0 );
    d_8 : in std_logic_vector( 1-1 downto 0 );
    d_9 : in std_logic_vector( 1-1 downto 0 );
    d_10 : in std_logic_vector( 1-1 downto 0 );
    d_11 : in std_logic_vector( 1-1 downto 0 );
    d_12 : in std_logic_vector( 1-1 downto 0 );
    d_13 : in std_logic_vector( 1-1 downto 0 );
    d_14 : in std_logic_vector( 1-1 downto 0 );
    d_15 : in std_logic_vector( 1-1 downto 0 );
    d_16 : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    q_1 : out std_logic_vector( 1-1 downto 0 );
    q_2 : out std_logic_vector( 1-1 downto 0 );
    q_3 : out std_logic_vector( 1-1 downto 0 );
    q_4 : out std_logic_vector( 1-1 downto 0 );
    q_5 : out std_logic_vector( 1-1 downto 0 );
    q_6 : out std_logic_vector( 1-1 downto 0 );
    q_7 : out std_logic_vector( 1-1 downto 0 );
    q_8 : out std_logic_vector( 1-1 downto 0 );
    q_9 : out std_logic_vector( 1-1 downto 0 );
    q_10 : out std_logic_vector( 1-1 downto 0 );
    q_11 : out std_logic_vector( 1-1 downto 0 );
    q_12 : out std_logic_vector( 1-1 downto 0 );
    q_13 : out std_logic_vector( 1-1 downto 0 );
    q_14 : out std_logic_vector( 1-1 downto 0 );
    q_15 : out std_logic_vector( 1-1 downto 0 );
    q_16 : out std_logic_vector( 1-1 downto 0 )
  );
end psb3_0_vector_delay1_x6;
architecture structural of psb3_0_vector_delay1_x6 is 
  signal delay0_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay12_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay9_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay15_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay10_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay13_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal ce_net : std_logic;
  signal slice3_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay14_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay7_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay11_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 1-1 downto 0 );
begin
  q_1 <= delay0_q_net;
  q_2 <= delay1_q_net;
  q_3 <= delay2_q_net;
  q_4 <= delay3_q_net;
  q_5 <= delay4_q_net;
  q_6 <= delay5_q_net;
  q_7 <= delay6_q_net;
  q_8 <= delay7_q_net;
  q_9 <= delay8_q_net;
  q_10 <= delay9_q_net;
  q_11 <= delay10_q_net;
  q_12 <= delay11_q_net;
  q_13 <= delay12_q_net;
  q_14 <= delay13_q_net;
  q_15 <= delay14_q_net;
  q_16 <= delay15_q_net;
  slice0_y_net <= d_1;
  slice1_y_net <= d_2;
  slice2_y_net <= d_3;
  slice3_y_net <= d_4;
  slice4_y_net <= d_5;
  slice5_y_net <= d_6;
  slice6_y_net <= d_7;
  slice7_y_net <= d_8;
  slice8_y_net <= d_9;
  slice9_y_net <= d_10;
  slice10_y_net <= d_11;
  slice11_y_net <= d_12;
  slice12_y_net <= d_13;
  slice13_y_net <= d_14;
  slice14_y_net <= d_15;
  slice15_y_net <= d_16;
  clk_net <= clk_1;
  ce_net <= ce_1;
  delay0 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice0_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay0_q_net
  );
  delay1 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice2_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay3 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice3_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  delay4 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice4_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net
  );
  delay5 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice5_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  delay6 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice6_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay6_q_net
  );
  delay7 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice7_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay7_q_net
  );
  delay8 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice8_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay8_q_net
  );
  delay9 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice9_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay9_q_net
  );
  delay10 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice10_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay10_q_net
  );
  delay11 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice11_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay11_q_net
  );
  delay12 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice12_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay12_q_net
  );
  delay13 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice13_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay13_q_net
  );
  delay14 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice14_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay14_q_net
  );
  delay15 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => slice15_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay15_q_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Overflow Detector add_re_4/Vector Slice
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_slice_x6 is
  port (
    in_1 : in std_logic_vector( 16-1 downto 0 );
    in_2 : in std_logic_vector( 16-1 downto 0 );
    in_3 : in std_logic_vector( 16-1 downto 0 );
    in_4 : in std_logic_vector( 16-1 downto 0 );
    in_5 : in std_logic_vector( 16-1 downto 0 );
    in_6 : in std_logic_vector( 16-1 downto 0 );
    in_7 : in std_logic_vector( 16-1 downto 0 );
    in_8 : in std_logic_vector( 16-1 downto 0 );
    in_9 : in std_logic_vector( 16-1 downto 0 );
    in_10 : in std_logic_vector( 16-1 downto 0 );
    in_11 : in std_logic_vector( 16-1 downto 0 );
    in_12 : in std_logic_vector( 16-1 downto 0 );
    in_13 : in std_logic_vector( 16-1 downto 0 );
    in_14 : in std_logic_vector( 16-1 downto 0 );
    in_15 : in std_logic_vector( 16-1 downto 0 );
    in_16 : in std_logic_vector( 16-1 downto 0 );
    out_1 : out std_logic_vector( 1-1 downto 0 );
    out_2 : out std_logic_vector( 1-1 downto 0 );
    out_3 : out std_logic_vector( 1-1 downto 0 );
    out_4 : out std_logic_vector( 1-1 downto 0 );
    out_5 : out std_logic_vector( 1-1 downto 0 );
    out_6 : out std_logic_vector( 1-1 downto 0 );
    out_7 : out std_logic_vector( 1-1 downto 0 );
    out_8 : out std_logic_vector( 1-1 downto 0 );
    out_9 : out std_logic_vector( 1-1 downto 0 );
    out_10 : out std_logic_vector( 1-1 downto 0 );
    out_11 : out std_logic_vector( 1-1 downto 0 );
    out_12 : out std_logic_vector( 1-1 downto 0 );
    out_13 : out std_logic_vector( 1-1 downto 0 );
    out_14 : out std_logic_vector( 1-1 downto 0 );
    out_15 : out std_logic_vector( 1-1 downto 0 );
    out_16 : out std_logic_vector( 1-1 downto 0 )
  );
end psb3_0_vector_slice_x6;
architecture structural of psb3_0_vector_slice_x6 is 
  signal slice10_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 1-1 downto 0 );
  signal mult0_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult1_p_net : std_logic_vector( 16-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 1-1 downto 0 );
  signal mult2_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult11_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult10_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult8_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult13_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult14_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult3_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult12_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult7_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult6_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult9_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult15_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult4_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult5_p_net : std_logic_vector( 16-1 downto 0 );
begin
  out_1 <= slice0_y_net;
  out_2 <= slice1_y_net;
  out_3 <= slice2_y_net;
  out_4 <= slice3_y_net;
  out_5 <= slice4_y_net;
  out_6 <= slice5_y_net;
  out_7 <= slice6_y_net;
  out_8 <= slice7_y_net;
  out_9 <= slice8_y_net;
  out_10 <= slice9_y_net;
  out_11 <= slice10_y_net;
  out_12 <= slice11_y_net;
  out_13 <= slice12_y_net;
  out_14 <= slice13_y_net;
  out_15 <= slice14_y_net;
  out_16 <= slice15_y_net;
  mult0_p_net <= in_1;
  mult1_p_net <= in_2;
  mult2_p_net <= in_3;
  mult3_p_net <= in_4;
  mult4_p_net <= in_5;
  mult5_p_net <= in_6;
  mult6_p_net <= in_7;
  mult7_p_net <= in_8;
  mult8_p_net <= in_9;
  mult9_p_net <= in_10;
  mult10_p_net <= in_11;
  mult11_p_net <= in_12;
  mult12_p_net <= in_13;
  mult13_p_net <= in_14;
  mult14_p_net <= in_15;
  mult15_p_net <= in_16;
  slice0 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult0_p_net,
    y => slice0_y_net
  );
  slice1 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult1_p_net,
    y => slice1_y_net
  );
  slice2 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult2_p_net,
    y => slice2_y_net
  );
  slice3 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult3_p_net,
    y => slice3_y_net
  );
  slice4 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult4_p_net,
    y => slice4_y_net
  );
  slice5 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult5_p_net,
    y => slice5_y_net
  );
  slice6 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult6_p_net,
    y => slice6_y_net
  );
  slice7 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult7_p_net,
    y => slice7_y_net
  );
  slice8 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult8_p_net,
    y => slice8_y_net
  );
  slice9 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult9_p_net,
    y => slice9_y_net
  );
  slice10 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult10_p_net,
    y => slice10_y_net
  );
  slice11 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult11_p_net,
    y => slice11_y_net
  );
  slice12 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult12_p_net,
    y => slice12_y_net
  );
  slice13 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult13_p_net,
    y => slice13_y_net
  );
  slice14 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult14_p_net,
    y => slice14_y_net
  );
  slice15 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => mult15_p_net,
    y => slice15_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Overflow Detector add_re_4/Vector Slice1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_slice1_x6 is
  port (
    in_1 : in std_logic_vector( 16-1 downto 0 );
    in_2 : in std_logic_vector( 16-1 downto 0 );
    in_3 : in std_logic_vector( 16-1 downto 0 );
    in_4 : in std_logic_vector( 16-1 downto 0 );
    in_5 : in std_logic_vector( 16-1 downto 0 );
    in_6 : in std_logic_vector( 16-1 downto 0 );
    in_7 : in std_logic_vector( 16-1 downto 0 );
    in_8 : in std_logic_vector( 16-1 downto 0 );
    in_9 : in std_logic_vector( 16-1 downto 0 );
    in_10 : in std_logic_vector( 16-1 downto 0 );
    in_11 : in std_logic_vector( 16-1 downto 0 );
    in_12 : in std_logic_vector( 16-1 downto 0 );
    in_13 : in std_logic_vector( 16-1 downto 0 );
    in_14 : in std_logic_vector( 16-1 downto 0 );
    in_15 : in std_logic_vector( 16-1 downto 0 );
    in_16 : in std_logic_vector( 16-1 downto 0 );
    out_1 : out std_logic_vector( 1-1 downto 0 );
    out_2 : out std_logic_vector( 1-1 downto 0 );
    out_3 : out std_logic_vector( 1-1 downto 0 );
    out_4 : out std_logic_vector( 1-1 downto 0 );
    out_5 : out std_logic_vector( 1-1 downto 0 );
    out_6 : out std_logic_vector( 1-1 downto 0 );
    out_7 : out std_logic_vector( 1-1 downto 0 );
    out_8 : out std_logic_vector( 1-1 downto 0 );
    out_9 : out std_logic_vector( 1-1 downto 0 );
    out_10 : out std_logic_vector( 1-1 downto 0 );
    out_11 : out std_logic_vector( 1-1 downto 0 );
    out_12 : out std_logic_vector( 1-1 downto 0 );
    out_13 : out std_logic_vector( 1-1 downto 0 );
    out_14 : out std_logic_vector( 1-1 downto 0 );
    out_15 : out std_logic_vector( 1-1 downto 0 );
    out_16 : out std_logic_vector( 1-1 downto 0 )
  );
end psb3_0_vector_slice1_x6;
architecture structural of psb3_0_vector_slice1_x6 is 
  signal slice0_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 1-1 downto 0 );
begin
  out_1 <= slice0_y_net;
  out_2 <= slice1_y_net;
  out_3 <= slice2_y_net;
  out_4 <= slice3_y_net;
  out_5 <= slice4_y_net;
  out_6 <= slice5_y_net;
  out_7 <= slice6_y_net;
  out_8 <= slice7_y_net;
  out_9 <= slice8_y_net;
  out_10 <= slice9_y_net;
  out_11 <= slice10_y_net;
  out_12 <= slice11_y_net;
  out_13 <= slice12_y_net;
  out_14 <= slice13_y_net;
  out_15 <= slice14_y_net;
  out_16 <= slice15_y_net;
  reinterpret0_output_port_net <= in_1;
  reinterpret1_output_port_net <= in_2;
  reinterpret2_output_port_net <= in_3;
  reinterpret3_output_port_net <= in_4;
  reinterpret4_output_port_net <= in_5;
  reinterpret5_output_port_net <= in_6;
  reinterpret6_output_port_net <= in_7;
  reinterpret7_output_port_net <= in_8;
  reinterpret8_output_port_net <= in_9;
  reinterpret9_output_port_net <= in_10;
  reinterpret10_output_port_net <= in_11;
  reinterpret11_output_port_net <= in_12;
  reinterpret12_output_port_net <= in_13;
  reinterpret13_output_port_net <= in_14;
  reinterpret14_output_port_net <= in_15;
  reinterpret15_output_port_net <= in_16;
  slice0 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret0_output_port_net,
    y => slice0_y_net
  );
  slice1 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret1_output_port_net,
    y => slice1_y_net
  );
  slice2 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret2_output_port_net,
    y => slice2_y_net
  );
  slice3 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret3_output_port_net,
    y => slice3_y_net
  );
  slice4 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret4_output_port_net,
    y => slice4_y_net
  );
  slice5 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret5_output_port_net,
    y => slice5_y_net
  );
  slice6 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret6_output_port_net,
    y => slice6_y_net
  );
  slice7 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret7_output_port_net,
    y => slice7_y_net
  );
  slice8 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret8_output_port_net,
    y => slice8_y_net
  );
  slice9 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret9_output_port_net,
    y => slice9_y_net
  );
  slice10 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret10_output_port_net,
    y => slice10_y_net
  );
  slice11 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret11_output_port_net,
    y => slice11_y_net
  );
  slice12 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret12_output_port_net,
    y => slice12_y_net
  );
  slice13 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret13_output_port_net,
    y => slice13_y_net
  );
  slice14 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret14_output_port_net,
    y => slice14_y_net
  );
  slice15 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => reinterpret15_output_port_net,
    y => slice15_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Overflow Detector add_re_4/Vector Slice2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_slice2_x6 is
  port (
    in_1 : in std_logic_vector( 16-1 downto 0 );
    in_2 : in std_logic_vector( 16-1 downto 0 );
    in_3 : in std_logic_vector( 16-1 downto 0 );
    in_4 : in std_logic_vector( 16-1 downto 0 );
    in_5 : in std_logic_vector( 16-1 downto 0 );
    in_6 : in std_logic_vector( 16-1 downto 0 );
    in_7 : in std_logic_vector( 16-1 downto 0 );
    in_8 : in std_logic_vector( 16-1 downto 0 );
    in_9 : in std_logic_vector( 16-1 downto 0 );
    in_10 : in std_logic_vector( 16-1 downto 0 );
    in_11 : in std_logic_vector( 16-1 downto 0 );
    in_12 : in std_logic_vector( 16-1 downto 0 );
    in_13 : in std_logic_vector( 16-1 downto 0 );
    in_14 : in std_logic_vector( 16-1 downto 0 );
    in_15 : in std_logic_vector( 16-1 downto 0 );
    in_16 : in std_logic_vector( 16-1 downto 0 );
    out_1 : out std_logic_vector( 1-1 downto 0 );
    out_2 : out std_logic_vector( 1-1 downto 0 );
    out_3 : out std_logic_vector( 1-1 downto 0 );
    out_4 : out std_logic_vector( 1-1 downto 0 );
    out_5 : out std_logic_vector( 1-1 downto 0 );
    out_6 : out std_logic_vector( 1-1 downto 0 );
    out_7 : out std_logic_vector( 1-1 downto 0 );
    out_8 : out std_logic_vector( 1-1 downto 0 );
    out_9 : out std_logic_vector( 1-1 downto 0 );
    out_10 : out std_logic_vector( 1-1 downto 0 );
    out_11 : out std_logic_vector( 1-1 downto 0 );
    out_12 : out std_logic_vector( 1-1 downto 0 );
    out_13 : out std_logic_vector( 1-1 downto 0 );
    out_14 : out std_logic_vector( 1-1 downto 0 );
    out_15 : out std_logic_vector( 1-1 downto 0 );
    out_16 : out std_logic_vector( 1-1 downto 0 )
  );
end psb3_0_vector_slice2_x6;
architecture structural of psb3_0_vector_slice2_x6 is 
  signal slice6_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 1-1 downto 0 );
  signal addsub0_s_net : std_logic_vector( 16-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 1-1 downto 0 );
  signal addsub13_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub9_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub6_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub12_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub3_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub7_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub11_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub14_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub8_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub5_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub10_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub15_s_net : std_logic_vector( 16-1 downto 0 );
begin
  out_1 <= slice0_y_net;
  out_2 <= slice1_y_net;
  out_3 <= slice2_y_net;
  out_4 <= slice3_y_net;
  out_5 <= slice4_y_net;
  out_6 <= slice5_y_net;
  out_7 <= slice6_y_net;
  out_8 <= slice7_y_net;
  out_9 <= slice8_y_net;
  out_10 <= slice9_y_net;
  out_11 <= slice10_y_net;
  out_12 <= slice11_y_net;
  out_13 <= slice12_y_net;
  out_14 <= slice13_y_net;
  out_15 <= slice14_y_net;
  out_16 <= slice15_y_net;
  addsub0_s_net <= in_1;
  addsub1_s_net <= in_2;
  addsub2_s_net <= in_3;
  addsub3_s_net <= in_4;
  addsub4_s_net <= in_5;
  addsub5_s_net <= in_6;
  addsub6_s_net <= in_7;
  addsub7_s_net <= in_8;
  addsub8_s_net <= in_9;
  addsub9_s_net <= in_10;
  addsub10_s_net <= in_11;
  addsub11_s_net <= in_12;
  addsub12_s_net <= in_13;
  addsub13_s_net <= in_14;
  addsub14_s_net <= in_15;
  addsub15_s_net <= in_16;
  slice0 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub0_s_net,
    y => slice0_y_net
  );
  slice1 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub1_s_net,
    y => slice1_y_net
  );
  slice2 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub2_s_net,
    y => slice2_y_net
  );
  slice3 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub3_s_net,
    y => slice3_y_net
  );
  slice4 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub4_s_net,
    y => slice4_y_net
  );
  slice5 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub5_s_net,
    y => slice5_y_net
  );
  slice6 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub6_s_net,
    y => slice6_y_net
  );
  slice7 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub7_s_net,
    y => slice7_y_net
  );
  slice8 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub8_s_net,
    y => slice8_y_net
  );
  slice9 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub9_s_net,
    y => slice9_y_net
  );
  slice10 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub10_s_net,
    y => slice10_y_net
  );
  slice11 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub11_s_net,
    y => slice11_y_net
  );
  slice12 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub12_s_net,
    y => slice12_y_net
  );
  slice13 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub13_s_net,
    y => slice13_y_net
  );
  slice14 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub14_s_net,
    y => slice14_y_net
  );
  slice15 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 15,
    new_msb => 15,
    x_width => 16,
    y_width => 1
  )
  port map (
    x => addsub15_s_net,
    y => slice15_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Overflow Detector add_re_4/Vector to Scalar
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_to_scalar_x6 is
  port (
    i_1 : in std_logic_vector( 1-1 downto 0 );
    i_2 : in std_logic_vector( 1-1 downto 0 );
    i_3 : in std_logic_vector( 1-1 downto 0 );
    i_4 : in std_logic_vector( 1-1 downto 0 );
    i_5 : in std_logic_vector( 1-1 downto 0 );
    i_6 : in std_logic_vector( 1-1 downto 0 );
    i_7 : in std_logic_vector( 1-1 downto 0 );
    i_8 : in std_logic_vector( 1-1 downto 0 );
    i_9 : in std_logic_vector( 1-1 downto 0 );
    i_10 : in std_logic_vector( 1-1 downto 0 );
    i_11 : in std_logic_vector( 1-1 downto 0 );
    i_12 : in std_logic_vector( 1-1 downto 0 );
    i_13 : in std_logic_vector( 1-1 downto 0 );
    i_14 : in std_logic_vector( 1-1 downto 0 );
    i_15 : in std_logic_vector( 1-1 downto 0 );
    i_16 : in std_logic_vector( 1-1 downto 0 );
    o : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_vector_to_scalar_x6;
architecture structural of psb3_0_vector_to_scalar_x6 is 
  signal concat1_y_net : std_logic_vector( 16-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay12_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay13_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay14_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay9_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay10_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay7_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay15_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay0_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay11_q_net : std_logic_vector( 1-1 downto 0 );
begin
  o <= concat1_y_net;
  delay0_q_net <= i_1;
  delay1_q_net <= i_2;
  delay2_q_net <= i_3;
  delay3_q_net <= i_4;
  delay4_q_net <= i_5;
  delay5_q_net <= i_6;
  delay6_q_net <= i_7;
  delay7_q_net <= i_8;
  delay8_q_net <= i_9;
  delay9_q_net <= i_10;
  delay10_q_net <= i_11;
  delay11_q_net <= i_12;
  delay12_q_net <= i_13;
  delay13_q_net <= i_14;
  delay14_q_net <= i_15;
  delay15_q_net <= i_16;
  concat1 : entity xil_defaultlib.sysgen_concat_d977c66e35 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => delay15_q_net,
    in1 => delay14_q_net,
    in2 => delay13_q_net,
    in3 => delay12_q_net,
    in4 => delay11_q_net,
    in5 => delay10_q_net,
    in6 => delay9_q_net,
    in7 => delay8_q_net,
    in8 => delay7_q_net,
    in9 => delay6_q_net,
    in10 => delay5_q_net,
    in11 => delay4_q_net,
    in12 => delay3_q_net,
    in13 => delay2_q_net,
    in14 => delay1_q_net,
    in15 => delay0_q_net,
    y => concat1_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Overflow Detector add_re_4/Vector to Scalar1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_to_scalar1_x6 is
  port (
    i_1 : in std_logic_vector( 1-1 downto 0 );
    i_2 : in std_logic_vector( 1-1 downto 0 );
    i_3 : in std_logic_vector( 1-1 downto 0 );
    i_4 : in std_logic_vector( 1-1 downto 0 );
    i_5 : in std_logic_vector( 1-1 downto 0 );
    i_6 : in std_logic_vector( 1-1 downto 0 );
    i_7 : in std_logic_vector( 1-1 downto 0 );
    i_8 : in std_logic_vector( 1-1 downto 0 );
    i_9 : in std_logic_vector( 1-1 downto 0 );
    i_10 : in std_logic_vector( 1-1 downto 0 );
    i_11 : in std_logic_vector( 1-1 downto 0 );
    i_12 : in std_logic_vector( 1-1 downto 0 );
    i_13 : in std_logic_vector( 1-1 downto 0 );
    i_14 : in std_logic_vector( 1-1 downto 0 );
    i_15 : in std_logic_vector( 1-1 downto 0 );
    i_16 : in std_logic_vector( 1-1 downto 0 );
    o : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_vector_to_scalar1_x6;
architecture structural of psb3_0_vector_to_scalar1_x6 is 
  signal delay14_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay11_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay12_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay10_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay15_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay9_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay7_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay13_q_net : std_logic_vector( 1-1 downto 0 );
  signal concat1_y_net : std_logic_vector( 16-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay0_q_net : std_logic_vector( 1-1 downto 0 );
begin
  o <= concat1_y_net;
  delay0_q_net <= i_1;
  delay1_q_net <= i_2;
  delay2_q_net <= i_3;
  delay3_q_net <= i_4;
  delay4_q_net <= i_5;
  delay5_q_net <= i_6;
  delay6_q_net <= i_7;
  delay7_q_net <= i_8;
  delay8_q_net <= i_9;
  delay9_q_net <= i_10;
  delay10_q_net <= i_11;
  delay11_q_net <= i_12;
  delay12_q_net <= i_13;
  delay13_q_net <= i_14;
  delay14_q_net <= i_15;
  delay15_q_net <= i_16;
  concat1 : entity xil_defaultlib.sysgen_concat_d977c66e35 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => delay15_q_net,
    in1 => delay14_q_net,
    in2 => delay13_q_net,
    in3 => delay12_q_net,
    in4 => delay11_q_net,
    in5 => delay10_q_net,
    in6 => delay9_q_net,
    in7 => delay8_q_net,
    in8 => delay7_q_net,
    in9 => delay6_q_net,
    in10 => delay5_q_net,
    in11 => delay4_q_net,
    in12 => delay3_q_net,
    in13 => delay2_q_net,
    in14 => delay1_q_net,
    in15 => delay0_q_net,
    y => concat1_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Overflow Detector add_re_4/Vector to Scalar2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_to_scalar2_x6 is
  port (
    i_1 : in std_logic_vector( 1-1 downto 0 );
    i_2 : in std_logic_vector( 1-1 downto 0 );
    i_3 : in std_logic_vector( 1-1 downto 0 );
    i_4 : in std_logic_vector( 1-1 downto 0 );
    i_5 : in std_logic_vector( 1-1 downto 0 );
    i_6 : in std_logic_vector( 1-1 downto 0 );
    i_7 : in std_logic_vector( 1-1 downto 0 );
    i_8 : in std_logic_vector( 1-1 downto 0 );
    i_9 : in std_logic_vector( 1-1 downto 0 );
    i_10 : in std_logic_vector( 1-1 downto 0 );
    i_11 : in std_logic_vector( 1-1 downto 0 );
    i_12 : in std_logic_vector( 1-1 downto 0 );
    i_13 : in std_logic_vector( 1-1 downto 0 );
    i_14 : in std_logic_vector( 1-1 downto 0 );
    i_15 : in std_logic_vector( 1-1 downto 0 );
    i_16 : in std_logic_vector( 1-1 downto 0 );
    o : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_vector_to_scalar2_x6;
architecture structural of psb3_0_vector_to_scalar2_x6 is 
  signal slice2_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 1-1 downto 0 );
  signal concat1_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 1-1 downto 0 );
begin
  o <= concat1_y_net;
  slice0_y_net <= i_1;
  slice1_y_net <= i_2;
  slice2_y_net <= i_3;
  slice3_y_net <= i_4;
  slice4_y_net <= i_5;
  slice5_y_net <= i_6;
  slice6_y_net <= i_7;
  slice7_y_net <= i_8;
  slice8_y_net <= i_9;
  slice9_y_net <= i_10;
  slice10_y_net <= i_11;
  slice11_y_net <= i_12;
  slice12_y_net <= i_13;
  slice13_y_net <= i_14;
  slice14_y_net <= i_15;
  slice15_y_net <= i_16;
  concat1 : entity xil_defaultlib.sysgen_concat_d977c66e35 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => slice15_y_net,
    in1 => slice14_y_net,
    in2 => slice13_y_net,
    in3 => slice12_y_net,
    in4 => slice11_y_net,
    in5 => slice10_y_net,
    in6 => slice9_y_net,
    in7 => slice8_y_net,
    in8 => slice7_y_net,
    in9 => slice6_y_net,
    in10 => slice5_y_net,
    in11 => slice4_y_net,
    in12 => slice3_y_net,
    in13 => slice2_y_net,
    in14 => slice1_y_net,
    in15 => slice0_y_net,
    y => concat1_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Overflow Detector add_re_4
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_overflow_detector_add_re_4 is
  port (
    rst : in std_logic_vector( 1-1 downto 0 );
    a_1 : in std_logic_vector( 16-1 downto 0 );
    b_1 : in std_logic_vector( 16-1 downto 0 );
    s_1 : in std_logic_vector( 16-1 downto 0 );
    a_2 : in std_logic_vector( 16-1 downto 0 );
    a_3 : in std_logic_vector( 16-1 downto 0 );
    a_4 : in std_logic_vector( 16-1 downto 0 );
    a_5 : in std_logic_vector( 16-1 downto 0 );
    a_6 : in std_logic_vector( 16-1 downto 0 );
    a_7 : in std_logic_vector( 16-1 downto 0 );
    a_8 : in std_logic_vector( 16-1 downto 0 );
    a_9 : in std_logic_vector( 16-1 downto 0 );
    a_10 : in std_logic_vector( 16-1 downto 0 );
    a_11 : in std_logic_vector( 16-1 downto 0 );
    a_12 : in std_logic_vector( 16-1 downto 0 );
    a_13 : in std_logic_vector( 16-1 downto 0 );
    a_14 : in std_logic_vector( 16-1 downto 0 );
    a_15 : in std_logic_vector( 16-1 downto 0 );
    a_16 : in std_logic_vector( 16-1 downto 0 );
    b_2 : in std_logic_vector( 16-1 downto 0 );
    b_3 : in std_logic_vector( 16-1 downto 0 );
    b_4 : in std_logic_vector( 16-1 downto 0 );
    b_5 : in std_logic_vector( 16-1 downto 0 );
    b_6 : in std_logic_vector( 16-1 downto 0 );
    b_7 : in std_logic_vector( 16-1 downto 0 );
    b_8 : in std_logic_vector( 16-1 downto 0 );
    b_9 : in std_logic_vector( 16-1 downto 0 );
    b_10 : in std_logic_vector( 16-1 downto 0 );
    b_11 : in std_logic_vector( 16-1 downto 0 );
    b_12 : in std_logic_vector( 16-1 downto 0 );
    b_13 : in std_logic_vector( 16-1 downto 0 );
    b_14 : in std_logic_vector( 16-1 downto 0 );
    b_15 : in std_logic_vector( 16-1 downto 0 );
    b_16 : in std_logic_vector( 16-1 downto 0 );
    s_2 : in std_logic_vector( 16-1 downto 0 );
    s_3 : in std_logic_vector( 16-1 downto 0 );
    s_4 : in std_logic_vector( 16-1 downto 0 );
    s_5 : in std_logic_vector( 16-1 downto 0 );
    s_6 : in std_logic_vector( 16-1 downto 0 );
    s_7 : in std_logic_vector( 16-1 downto 0 );
    s_8 : in std_logic_vector( 16-1 downto 0 );
    s_9 : in std_logic_vector( 16-1 downto 0 );
    s_10 : in std_logic_vector( 16-1 downto 0 );
    s_11 : in std_logic_vector( 16-1 downto 0 );
    s_12 : in std_logic_vector( 16-1 downto 0 );
    s_13 : in std_logic_vector( 16-1 downto 0 );
    s_14 : in std_logic_vector( 16-1 downto 0 );
    s_15 : in std_logic_vector( 16-1 downto 0 );
    s_16 : in std_logic_vector( 16-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    ov : out std_logic_vector( 1-1 downto 0 )
  );
end psb3_0_overflow_detector_add_re_4;
architecture structural of psb3_0_overflow_detector_add_re_4 is 
  signal mult1_p_net : std_logic_vector( 16-1 downto 0 );
  signal gin_tl_reset_net : std_logic_vector( 1-1 downto 0 );
  signal mult5_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult6_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult7_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult8_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mult2_p_net : std_logic_vector( 16-1 downto 0 );
  signal register_q_net : std_logic_vector( 1-1 downto 0 );
  signal mult0_p_net : std_logic_vector( 16-1 downto 0 );
  signal addsub0_s_net : std_logic_vector( 16-1 downto 0 );
  signal mult3_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult4_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult9_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub3_s_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 16-1 downto 0 );
  signal mult15_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mult12_p_net : std_logic_vector( 16-1 downto 0 );
  signal addsub7_s_net : std_logic_vector( 16-1 downto 0 );
  signal mult11_p_net : std_logic_vector( 16-1 downto 0 );
  signal addsub8_s_net : std_logic_vector( 16-1 downto 0 );
  signal mult10_p_net : std_logic_vector( 16-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub5_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub6_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub9_s_net : std_logic_vector( 16-1 downto 0 );
  signal mult13_p_net : std_logic_vector( 16-1 downto 0 );
  signal addsub10_s_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mult14_p_net : std_logic_vector( 16-1 downto 0 );
  signal slice0_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal slice4_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal slice13_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 1-1 downto 0 );
  signal addsub13_s_net : std_logic_vector( 16-1 downto 0 );
  signal slice5_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal slice7_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal delay5_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay6_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice11_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal delay0_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay14_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal slice15_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay11_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay15_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal addsub15_s_net : std_logic_vector( 16-1 downto 0 );
  signal delay0_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice2_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal slice8_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal slice6_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal slice9_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal delay12_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay10_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal addsub12_s_net : std_logic_vector( 16-1 downto 0 );
  signal delay4_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay7_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice12_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice1_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal delay8_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice3_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal addsub14_s_net : std_logic_vector( 16-1 downto 0 );
  signal delay1_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay9_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay13_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay13_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay10_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay14_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay11_q_net : std_logic_vector( 1-1 downto 0 );
  signal addsub11_s_net : std_logic_vector( 16-1 downto 0 );
  signal delay3_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay7_q_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal slice10_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal delay12_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay15_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice0_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice1_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice2_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice14_y_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal delay9_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice5_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice3_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice11_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice12_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 1-1 downto 0 );
  signal concat1_y_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal concat1_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 1-1 downto 0 );
  signal concat1_y_net_x1 : std_logic_vector( 16-1 downto 0 );
  signal slice6_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice7_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice9_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice15_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal expression_dout_net : std_logic_vector( 1-1 downto 0 );
  signal slice8_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 1-1 downto 0 );
  signal constant17_op_net : std_logic_vector( 1-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 1-1 downto 0 );
  signal convert_dout_net : std_logic_vector( 1-1 downto 0 );
  signal slice10_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice4_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice14_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice13_y_net_x0 : std_logic_vector( 1-1 downto 0 );
begin
  ov <= register_q_net;
  gin_tl_reset_net <= rst;
  mult0_p_net <= a_1;
  reinterpret0_output_port_net <= b_1;
  addsub0_s_net <= s_1;
  mult1_p_net <= a_2;
  mult2_p_net <= a_3;
  mult3_p_net <= a_4;
  mult4_p_net <= a_5;
  mult5_p_net <= a_6;
  mult6_p_net <= a_7;
  mult7_p_net <= a_8;
  mult8_p_net <= a_9;
  mult9_p_net <= a_10;
  mult10_p_net <= a_11;
  mult11_p_net <= a_12;
  mult12_p_net <= a_13;
  mult13_p_net <= a_14;
  mult14_p_net <= a_15;
  mult15_p_net <= a_16;
  reinterpret1_output_port_net <= b_2;
  reinterpret2_output_port_net <= b_3;
  reinterpret3_output_port_net <= b_4;
  reinterpret4_output_port_net <= b_5;
  reinterpret5_output_port_net <= b_6;
  reinterpret6_output_port_net <= b_7;
  reinterpret7_output_port_net <= b_8;
  reinterpret8_output_port_net <= b_9;
  reinterpret9_output_port_net <= b_10;
  reinterpret10_output_port_net <= b_11;
  reinterpret11_output_port_net <= b_12;
  reinterpret12_output_port_net <= b_13;
  reinterpret13_output_port_net <= b_14;
  reinterpret14_output_port_net <= b_15;
  reinterpret15_output_port_net <= b_16;
  addsub1_s_net <= s_2;
  addsub2_s_net <= s_3;
  addsub3_s_net <= s_4;
  addsub4_s_net <= s_5;
  addsub5_s_net <= s_6;
  addsub6_s_net <= s_7;
  addsub7_s_net <= s_8;
  addsub8_s_net <= s_9;
  addsub9_s_net <= s_10;
  addsub10_s_net <= s_11;
  addsub11_s_net <= s_12;
  addsub12_s_net <= s_13;
  addsub13_s_net <= s_14;
  addsub14_s_net <= s_15;
  addsub15_s_net <= s_16;
  clk_net <= clk_1;
  ce_net <= ce_1;
  vector_delay : entity xil_defaultlib.psb3_0_vector_delay_x6 
  port map (
    d_1 => slice0_y_net_x1,
    d_2 => slice1_y_net_x1,
    d_3 => slice2_y_net_x1,
    d_4 => slice3_y_net_x1,
    d_5 => slice4_y_net_x1,
    d_6 => slice5_y_net_x1,
    d_7 => slice6_y_net_x1,
    d_8 => slice7_y_net_x1,
    d_9 => slice8_y_net_x1,
    d_10 => slice9_y_net_x1,
    d_11 => slice10_y_net_x1,
    d_12 => slice11_y_net_x1,
    d_13 => slice12_y_net_x1,
    d_14 => slice13_y_net_x1,
    d_15 => slice14_y_net_x1,
    d_16 => slice15_y_net_x1,
    clk_1 => clk_net,
    ce_1 => ce_net,
    q_1 => delay0_q_net_x0,
    q_2 => delay1_q_net_x0,
    q_3 => delay2_q_net_x0,
    q_4 => delay3_q_net_x0,
    q_5 => delay4_q_net_x0,
    q_6 => delay5_q_net_x0,
    q_7 => delay6_q_net_x0,
    q_8 => delay7_q_net_x0,
    q_9 => delay8_q_net_x0,
    q_10 => delay9_q_net_x0,
    q_11 => delay10_q_net_x0,
    q_12 => delay11_q_net_x0,
    q_13 => delay12_q_net_x0,
    q_14 => delay13_q_net_x0,
    q_15 => delay14_q_net_x0,
    q_16 => delay15_q_net_x0
  );
  vector_delay1 : entity xil_defaultlib.psb3_0_vector_delay1_x6 
  port map (
    d_1 => slice0_y_net_x0,
    d_2 => slice1_y_net_x0,
    d_3 => slice2_y_net_x0,
    d_4 => slice3_y_net_x0,
    d_5 => slice4_y_net_x0,
    d_6 => slice5_y_net_x0,
    d_7 => slice6_y_net_x0,
    d_8 => slice7_y_net_x0,
    d_9 => slice8_y_net_x0,
    d_10 => slice9_y_net_x0,
    d_11 => slice10_y_net_x0,
    d_12 => slice11_y_net_x0,
    d_13 => slice12_y_net_x0,
    d_14 => slice13_y_net_x0,
    d_15 => slice14_y_net_x0,
    d_16 => slice15_y_net_x0,
    clk_1 => clk_net,
    ce_1 => ce_net,
    q_1 => delay0_q_net,
    q_2 => delay1_q_net,
    q_3 => delay2_q_net,
    q_4 => delay3_q_net,
    q_5 => delay4_q_net,
    q_6 => delay5_q_net,
    q_7 => delay6_q_net,
    q_8 => delay7_q_net,
    q_9 => delay8_q_net,
    q_10 => delay9_q_net,
    q_11 => delay10_q_net,
    q_12 => delay11_q_net,
    q_13 => delay12_q_net,
    q_14 => delay13_q_net,
    q_15 => delay14_q_net,
    q_16 => delay15_q_net
  );
  vector_slice : entity xil_defaultlib.psb3_0_vector_slice_x6 
  port map (
    in_1 => mult0_p_net,
    in_2 => mult1_p_net,
    in_3 => mult2_p_net,
    in_4 => mult3_p_net,
    in_5 => mult4_p_net,
    in_6 => mult5_p_net,
    in_7 => mult6_p_net,
    in_8 => mult7_p_net,
    in_9 => mult8_p_net,
    in_10 => mult9_p_net,
    in_11 => mult10_p_net,
    in_12 => mult11_p_net,
    in_13 => mult12_p_net,
    in_14 => mult13_p_net,
    in_15 => mult14_p_net,
    in_16 => mult15_p_net,
    out_1 => slice0_y_net_x1,
    out_2 => slice1_y_net_x1,
    out_3 => slice2_y_net_x1,
    out_4 => slice3_y_net_x1,
    out_5 => slice4_y_net_x1,
    out_6 => slice5_y_net_x1,
    out_7 => slice6_y_net_x1,
    out_8 => slice7_y_net_x1,
    out_9 => slice8_y_net_x1,
    out_10 => slice9_y_net_x1,
    out_11 => slice10_y_net_x1,
    out_12 => slice11_y_net_x1,
    out_13 => slice12_y_net_x1,
    out_14 => slice13_y_net_x1,
    out_15 => slice14_y_net_x1,
    out_16 => slice15_y_net_x1
  );
  vector_slice1 : entity xil_defaultlib.psb3_0_vector_slice1_x6 
  port map (
    in_1 => reinterpret0_output_port_net,
    in_2 => reinterpret1_output_port_net,
    in_3 => reinterpret2_output_port_net,
    in_4 => reinterpret3_output_port_net,
    in_5 => reinterpret4_output_port_net,
    in_6 => reinterpret5_output_port_net,
    in_7 => reinterpret6_output_port_net,
    in_8 => reinterpret7_output_port_net,
    in_9 => reinterpret8_output_port_net,
    in_10 => reinterpret9_output_port_net,
    in_11 => reinterpret10_output_port_net,
    in_12 => reinterpret11_output_port_net,
    in_13 => reinterpret12_output_port_net,
    in_14 => reinterpret13_output_port_net,
    in_15 => reinterpret14_output_port_net,
    in_16 => reinterpret15_output_port_net,
    out_1 => slice0_y_net_x0,
    out_2 => slice1_y_net_x0,
    out_3 => slice2_y_net_x0,
    out_4 => slice3_y_net_x0,
    out_5 => slice4_y_net_x0,
    out_6 => slice5_y_net_x0,
    out_7 => slice6_y_net_x0,
    out_8 => slice7_y_net_x0,
    out_9 => slice8_y_net_x0,
    out_10 => slice9_y_net_x0,
    out_11 => slice10_y_net_x0,
    out_12 => slice11_y_net_x0,
    out_13 => slice12_y_net_x0,
    out_14 => slice13_y_net_x0,
    out_15 => slice14_y_net_x0,
    out_16 => slice15_y_net_x0
  );
  vector_slice2 : entity xil_defaultlib.psb3_0_vector_slice2_x6 
  port map (
    in_1 => addsub0_s_net,
    in_2 => addsub1_s_net,
    in_3 => addsub2_s_net,
    in_4 => addsub3_s_net,
    in_5 => addsub4_s_net,
    in_6 => addsub5_s_net,
    in_7 => addsub6_s_net,
    in_8 => addsub7_s_net,
    in_9 => addsub8_s_net,
    in_10 => addsub9_s_net,
    in_11 => addsub10_s_net,
    in_12 => addsub11_s_net,
    in_13 => addsub12_s_net,
    in_14 => addsub13_s_net,
    in_15 => addsub14_s_net,
    in_16 => addsub15_s_net,
    out_1 => slice0_y_net,
    out_2 => slice1_y_net,
    out_3 => slice2_y_net,
    out_4 => slice3_y_net,
    out_5 => slice4_y_net,
    out_6 => slice5_y_net,
    out_7 => slice6_y_net,
    out_8 => slice7_y_net,
    out_9 => slice8_y_net,
    out_10 => slice9_y_net,
    out_11 => slice10_y_net,
    out_12 => slice11_y_net,
    out_13 => slice12_y_net,
    out_14 => slice13_y_net,
    out_15 => slice14_y_net,
    out_16 => slice15_y_net
  );
  vector_to_scalar : entity xil_defaultlib.psb3_0_vector_to_scalar_x6 
  port map (
    i_1 => delay0_q_net_x0,
    i_2 => delay1_q_net_x0,
    i_3 => delay2_q_net_x0,
    i_4 => delay3_q_net_x0,
    i_5 => delay4_q_net_x0,
    i_6 => delay5_q_net_x0,
    i_7 => delay6_q_net_x0,
    i_8 => delay7_q_net_x0,
    i_9 => delay8_q_net_x0,
    i_10 => delay9_q_net_x0,
    i_11 => delay10_q_net_x0,
    i_12 => delay11_q_net_x0,
    i_13 => delay12_q_net_x0,
    i_14 => delay13_q_net_x0,
    i_15 => delay14_q_net_x0,
    i_16 => delay15_q_net_x0,
    o => concat1_y_net_x1
  );
  vector_to_scalar1 : entity xil_defaultlib.psb3_0_vector_to_scalar1_x6 
  port map (
    i_1 => delay0_q_net,
    i_2 => delay1_q_net,
    i_3 => delay2_q_net,
    i_4 => delay3_q_net,
    i_5 => delay4_q_net,
    i_6 => delay5_q_net,
    i_7 => delay6_q_net,
    i_8 => delay7_q_net,
    i_9 => delay8_q_net,
    i_10 => delay9_q_net,
    i_11 => delay10_q_net,
    i_12 => delay11_q_net,
    i_13 => delay12_q_net,
    i_14 => delay13_q_net,
    i_15 => delay14_q_net,
    i_16 => delay15_q_net,
    o => concat1_y_net_x0
  );
  vector_to_scalar2 : entity xil_defaultlib.psb3_0_vector_to_scalar2_x6 
  port map (
    i_1 => slice0_y_net,
    i_2 => slice1_y_net,
    i_3 => slice2_y_net,
    i_4 => slice3_y_net,
    i_5 => slice4_y_net,
    i_6 => slice5_y_net,
    i_7 => slice6_y_net,
    i_8 => slice7_y_net,
    i_9 => slice8_y_net,
    i_10 => slice9_y_net,
    i_11 => slice10_y_net,
    i_12 => slice11_y_net,
    i_13 => slice12_y_net,
    i_14 => slice13_y_net,
    i_15 => slice14_y_net,
    i_16 => slice15_y_net,
    o => concat1_y_net
  );
  constant17 : entity xil_defaultlib.sysgen_constant_71e89d757c 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant17_op_net
  );
  convert : entity xil_defaultlib.psb3_0_xlconvert 
  generic map (
    bool_conversion => 1,
    din_arith => 1,
    din_bin_pt => 0,
    din_width => 1,
    dout_arith => 1,
    dout_bin_pt => 0,
    dout_width => 1,
    latency => 1,
    overflow => xlWrap,
    quantization => xlTruncate
  )
  port map (
    clr => '0',
    en => "1",
    din => expression_dout_net,
    clk => clk_net,
    ce => ce_net,
    dout => convert_dout_net
  );
  expression : entity xil_defaultlib.sysgen_expr_7c83532765 
  port map (
    clr => '0',
    a => concat1_y_net_x1,
    b => concat1_y_net_x0,
    s => concat1_y_net,
    clk => clk_net,
    ce => ce_net,
    dout => expression_dout_net
  );
  register_x0 : entity xil_defaultlib.psb3_0_xlregister 
  generic map (
    d_width => 1,
    init_value => b"0"
  )
  port map (
    d => constant17_op_net,
    rst => gin_tl_reset_net,
    en => convert_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => register_q_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Scalar to Vector1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_scalar_to_vector1 is
  port (
    i : in std_logic_vector( 256-1 downto 0 );
    o_1 : out std_logic_vector( 16-1 downto 0 );
    o_2 : out std_logic_vector( 16-1 downto 0 );
    o_3 : out std_logic_vector( 16-1 downto 0 );
    o_4 : out std_logic_vector( 16-1 downto 0 );
    o_5 : out std_logic_vector( 16-1 downto 0 );
    o_6 : out std_logic_vector( 16-1 downto 0 );
    o_7 : out std_logic_vector( 16-1 downto 0 );
    o_8 : out std_logic_vector( 16-1 downto 0 );
    o_9 : out std_logic_vector( 16-1 downto 0 );
    o_10 : out std_logic_vector( 16-1 downto 0 );
    o_11 : out std_logic_vector( 16-1 downto 0 );
    o_12 : out std_logic_vector( 16-1 downto 0 );
    o_13 : out std_logic_vector( 16-1 downto 0 );
    o_14 : out std_logic_vector( 16-1 downto 0 );
    o_15 : out std_logic_vector( 16-1 downto 0 );
    o_16 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_scalar_to_vector1;
architecture structural of psb3_0_scalar_to_vector1 is 
  signal slice1_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 16-1 downto 0 );
  signal bitbasher1_a_net : std_logic_vector( 256-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 16-1 downto 0 );
begin
  o_1 <= slice0_y_net;
  o_2 <= slice1_y_net;
  o_3 <= slice2_y_net;
  o_4 <= slice3_y_net;
  o_5 <= slice4_y_net;
  o_6 <= slice5_y_net;
  o_7 <= slice6_y_net;
  o_8 <= slice7_y_net;
  o_9 <= slice8_y_net;
  o_10 <= slice9_y_net;
  o_11 <= slice10_y_net;
  o_12 <= slice11_y_net;
  o_13 <= slice12_y_net;
  o_14 <= slice13_y_net;
  o_15 <= slice14_y_net;
  o_16 <= slice15_y_net;
  bitbasher1_a_net <= i;
  slice0 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 15,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher1_a_net,
    y => slice0_y_net
  );
  slice1 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 16,
    new_msb => 31,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher1_a_net,
    y => slice1_y_net
  );
  slice2 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 32,
    new_msb => 47,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher1_a_net,
    y => slice2_y_net
  );
  slice3 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 48,
    new_msb => 63,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher1_a_net,
    y => slice3_y_net
  );
  slice4 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 64,
    new_msb => 79,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher1_a_net,
    y => slice4_y_net
  );
  slice5 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 80,
    new_msb => 95,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher1_a_net,
    y => slice5_y_net
  );
  slice6 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 96,
    new_msb => 111,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher1_a_net,
    y => slice6_y_net
  );
  slice7 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 112,
    new_msb => 127,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher1_a_net,
    y => slice7_y_net
  );
  slice8 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 128,
    new_msb => 143,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher1_a_net,
    y => slice8_y_net
  );
  slice9 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 144,
    new_msb => 159,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher1_a_net,
    y => slice9_y_net
  );
  slice10 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 160,
    new_msb => 175,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher1_a_net,
    y => slice10_y_net
  );
  slice11 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 176,
    new_msb => 191,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher1_a_net,
    y => slice11_y_net
  );
  slice12 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 192,
    new_msb => 207,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher1_a_net,
    y => slice12_y_net
  );
  slice13 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 208,
    new_msb => 223,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher1_a_net,
    y => slice13_y_net
  );
  slice14 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 224,
    new_msb => 239,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher1_a_net,
    y => slice14_y_net
  );
  slice15 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 240,
    new_msb => 255,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher1_a_net,
    y => slice15_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Scalar to Vector2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_scalar_to_vector2 is
  port (
    i : in std_logic_vector( 256-1 downto 0 );
    o_1 : out std_logic_vector( 16-1 downto 0 );
    o_2 : out std_logic_vector( 16-1 downto 0 );
    o_3 : out std_logic_vector( 16-1 downto 0 );
    o_4 : out std_logic_vector( 16-1 downto 0 );
    o_5 : out std_logic_vector( 16-1 downto 0 );
    o_6 : out std_logic_vector( 16-1 downto 0 );
    o_7 : out std_logic_vector( 16-1 downto 0 );
    o_8 : out std_logic_vector( 16-1 downto 0 );
    o_9 : out std_logic_vector( 16-1 downto 0 );
    o_10 : out std_logic_vector( 16-1 downto 0 );
    o_11 : out std_logic_vector( 16-1 downto 0 );
    o_12 : out std_logic_vector( 16-1 downto 0 );
    o_13 : out std_logic_vector( 16-1 downto 0 );
    o_14 : out std_logic_vector( 16-1 downto 0 );
    o_15 : out std_logic_vector( 16-1 downto 0 );
    o_16 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_scalar_to_vector2;
architecture structural of psb3_0_scalar_to_vector2 is 
  signal slice0_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 16-1 downto 0 );
  signal bitbasher2_a_net : std_logic_vector( 256-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 16-1 downto 0 );
begin
  o_1 <= slice0_y_net;
  o_2 <= slice1_y_net;
  o_3 <= slice2_y_net;
  o_4 <= slice3_y_net;
  o_5 <= slice4_y_net;
  o_6 <= slice5_y_net;
  o_7 <= slice6_y_net;
  o_8 <= slice7_y_net;
  o_9 <= slice8_y_net;
  o_10 <= slice9_y_net;
  o_11 <= slice10_y_net;
  o_12 <= slice11_y_net;
  o_13 <= slice12_y_net;
  o_14 <= slice13_y_net;
  o_15 <= slice14_y_net;
  o_16 <= slice15_y_net;
  bitbasher2_a_net <= i;
  slice0 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 15,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher2_a_net,
    y => slice0_y_net
  );
  slice1 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 16,
    new_msb => 31,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher2_a_net,
    y => slice1_y_net
  );
  slice2 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 32,
    new_msb => 47,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher2_a_net,
    y => slice2_y_net
  );
  slice3 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 48,
    new_msb => 63,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher2_a_net,
    y => slice3_y_net
  );
  slice4 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 64,
    new_msb => 79,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher2_a_net,
    y => slice4_y_net
  );
  slice5 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 80,
    new_msb => 95,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher2_a_net,
    y => slice5_y_net
  );
  slice6 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 96,
    new_msb => 111,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher2_a_net,
    y => slice6_y_net
  );
  slice7 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 112,
    new_msb => 127,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher2_a_net,
    y => slice7_y_net
  );
  slice8 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 128,
    new_msb => 143,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher2_a_net,
    y => slice8_y_net
  );
  slice9 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 144,
    new_msb => 159,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher2_a_net,
    y => slice9_y_net
  );
  slice10 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 160,
    new_msb => 175,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher2_a_net,
    y => slice10_y_net
  );
  slice11 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 176,
    new_msb => 191,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher2_a_net,
    y => slice11_y_net
  );
  slice12 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 192,
    new_msb => 207,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher2_a_net,
    y => slice12_y_net
  );
  slice13 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 208,
    new_msb => 223,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher2_a_net,
    y => slice13_y_net
  );
  slice14 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 224,
    new_msb => 239,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher2_a_net,
    y => slice14_y_net
  );
  slice15 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 240,
    new_msb => 255,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher2_a_net,
    y => slice15_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Scalar to Vector3
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_scalar_to_vector3 is
  port (
    i : in std_logic_vector( 256-1 downto 0 );
    o_1 : out std_logic_vector( 16-1 downto 0 );
    o_2 : out std_logic_vector( 16-1 downto 0 );
    o_3 : out std_logic_vector( 16-1 downto 0 );
    o_4 : out std_logic_vector( 16-1 downto 0 );
    o_5 : out std_logic_vector( 16-1 downto 0 );
    o_6 : out std_logic_vector( 16-1 downto 0 );
    o_7 : out std_logic_vector( 16-1 downto 0 );
    o_8 : out std_logic_vector( 16-1 downto 0 );
    o_9 : out std_logic_vector( 16-1 downto 0 );
    o_10 : out std_logic_vector( 16-1 downto 0 );
    o_11 : out std_logic_vector( 16-1 downto 0 );
    o_12 : out std_logic_vector( 16-1 downto 0 );
    o_13 : out std_logic_vector( 16-1 downto 0 );
    o_14 : out std_logic_vector( 16-1 downto 0 );
    o_15 : out std_logic_vector( 16-1 downto 0 );
    o_16 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_scalar_to_vector3;
architecture structural of psb3_0_scalar_to_vector3 is 
  signal slice4_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 16-1 downto 0 );
  signal bitbasher3_a_net : std_logic_vector( 256-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 16-1 downto 0 );
begin
  o_1 <= slice0_y_net;
  o_2 <= slice1_y_net;
  o_3 <= slice2_y_net;
  o_4 <= slice3_y_net;
  o_5 <= slice4_y_net;
  o_6 <= slice5_y_net;
  o_7 <= slice6_y_net;
  o_8 <= slice7_y_net;
  o_9 <= slice8_y_net;
  o_10 <= slice9_y_net;
  o_11 <= slice10_y_net;
  o_12 <= slice11_y_net;
  o_13 <= slice12_y_net;
  o_14 <= slice13_y_net;
  o_15 <= slice14_y_net;
  o_16 <= slice15_y_net;
  bitbasher3_a_net <= i;
  slice0 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 15,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher3_a_net,
    y => slice0_y_net
  );
  slice1 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 16,
    new_msb => 31,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher3_a_net,
    y => slice1_y_net
  );
  slice2 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 32,
    new_msb => 47,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher3_a_net,
    y => slice2_y_net
  );
  slice3 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 48,
    new_msb => 63,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher3_a_net,
    y => slice3_y_net
  );
  slice4 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 64,
    new_msb => 79,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher3_a_net,
    y => slice4_y_net
  );
  slice5 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 80,
    new_msb => 95,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher3_a_net,
    y => slice5_y_net
  );
  slice6 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 96,
    new_msb => 111,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher3_a_net,
    y => slice6_y_net
  );
  slice7 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 112,
    new_msb => 127,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher3_a_net,
    y => slice7_y_net
  );
  slice8 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 128,
    new_msb => 143,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher3_a_net,
    y => slice8_y_net
  );
  slice9 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 144,
    new_msb => 159,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher3_a_net,
    y => slice9_y_net
  );
  slice10 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 160,
    new_msb => 175,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher3_a_net,
    y => slice10_y_net
  );
  slice11 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 176,
    new_msb => 191,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher3_a_net,
    y => slice11_y_net
  );
  slice12 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 192,
    new_msb => 207,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher3_a_net,
    y => slice12_y_net
  );
  slice13 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 208,
    new_msb => 223,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher3_a_net,
    y => slice13_y_net
  );
  slice14 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 224,
    new_msb => 239,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher3_a_net,
    y => slice14_y_net
  );
  slice15 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 240,
    new_msb => 255,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher3_a_net,
    y => slice15_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Scalar to Vector4
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_scalar_to_vector4 is
  port (
    i : in std_logic_vector( 256-1 downto 0 );
    o_1 : out std_logic_vector( 16-1 downto 0 );
    o_2 : out std_logic_vector( 16-1 downto 0 );
    o_3 : out std_logic_vector( 16-1 downto 0 );
    o_4 : out std_logic_vector( 16-1 downto 0 );
    o_5 : out std_logic_vector( 16-1 downto 0 );
    o_6 : out std_logic_vector( 16-1 downto 0 );
    o_7 : out std_logic_vector( 16-1 downto 0 );
    o_8 : out std_logic_vector( 16-1 downto 0 );
    o_9 : out std_logic_vector( 16-1 downto 0 );
    o_10 : out std_logic_vector( 16-1 downto 0 );
    o_11 : out std_logic_vector( 16-1 downto 0 );
    o_12 : out std_logic_vector( 16-1 downto 0 );
    o_13 : out std_logic_vector( 16-1 downto 0 );
    o_14 : out std_logic_vector( 16-1 downto 0 );
    o_15 : out std_logic_vector( 16-1 downto 0 );
    o_16 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_scalar_to_vector4;
architecture structural of psb3_0_scalar_to_vector4 is 
  signal slice6_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 16-1 downto 0 );
  signal bitbasher4_a_net : std_logic_vector( 256-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 16-1 downto 0 );
begin
  o_1 <= slice0_y_net;
  o_2 <= slice1_y_net;
  o_3 <= slice2_y_net;
  o_4 <= slice3_y_net;
  o_5 <= slice4_y_net;
  o_6 <= slice5_y_net;
  o_7 <= slice6_y_net;
  o_8 <= slice7_y_net;
  o_9 <= slice8_y_net;
  o_10 <= slice9_y_net;
  o_11 <= slice10_y_net;
  o_12 <= slice11_y_net;
  o_13 <= slice12_y_net;
  o_14 <= slice13_y_net;
  o_15 <= slice14_y_net;
  o_16 <= slice15_y_net;
  bitbasher4_a_net <= i;
  slice0 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 15,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher4_a_net,
    y => slice0_y_net
  );
  slice1 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 16,
    new_msb => 31,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher4_a_net,
    y => slice1_y_net
  );
  slice2 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 32,
    new_msb => 47,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher4_a_net,
    y => slice2_y_net
  );
  slice3 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 48,
    new_msb => 63,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher4_a_net,
    y => slice3_y_net
  );
  slice4 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 64,
    new_msb => 79,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher4_a_net,
    y => slice4_y_net
  );
  slice5 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 80,
    new_msb => 95,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher4_a_net,
    y => slice5_y_net
  );
  slice6 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 96,
    new_msb => 111,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher4_a_net,
    y => slice6_y_net
  );
  slice7 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 112,
    new_msb => 127,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher4_a_net,
    y => slice7_y_net
  );
  slice8 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 128,
    new_msb => 143,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher4_a_net,
    y => slice8_y_net
  );
  slice9 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 144,
    new_msb => 159,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher4_a_net,
    y => slice9_y_net
  );
  slice10 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 160,
    new_msb => 175,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher4_a_net,
    y => slice10_y_net
  );
  slice11 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 176,
    new_msb => 191,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher4_a_net,
    y => slice11_y_net
  );
  slice12 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 192,
    new_msb => 207,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher4_a_net,
    y => slice12_y_net
  );
  slice13 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 208,
    new_msb => 223,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher4_a_net,
    y => slice13_y_net
  );
  slice14 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 224,
    new_msb => 239,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher4_a_net,
    y => slice14_y_net
  );
  slice15 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 240,
    new_msb => 255,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher4_a_net,
    y => slice15_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Scalar to Vector5
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_scalar_to_vector5 is
  port (
    i : in std_logic_vector( 256-1 downto 0 );
    o_1 : out std_logic_vector( 16-1 downto 0 );
    o_2 : out std_logic_vector( 16-1 downto 0 );
    o_3 : out std_logic_vector( 16-1 downto 0 );
    o_4 : out std_logic_vector( 16-1 downto 0 );
    o_5 : out std_logic_vector( 16-1 downto 0 );
    o_6 : out std_logic_vector( 16-1 downto 0 );
    o_7 : out std_logic_vector( 16-1 downto 0 );
    o_8 : out std_logic_vector( 16-1 downto 0 );
    o_9 : out std_logic_vector( 16-1 downto 0 );
    o_10 : out std_logic_vector( 16-1 downto 0 );
    o_11 : out std_logic_vector( 16-1 downto 0 );
    o_12 : out std_logic_vector( 16-1 downto 0 );
    o_13 : out std_logic_vector( 16-1 downto 0 );
    o_14 : out std_logic_vector( 16-1 downto 0 );
    o_15 : out std_logic_vector( 16-1 downto 0 );
    o_16 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_scalar_to_vector5;
architecture structural of psb3_0_scalar_to_vector5 is 
  signal slice0_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 16-1 downto 0 );
  signal bitbasher5_a_net : std_logic_vector( 256-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 16-1 downto 0 );
begin
  o_1 <= slice0_y_net;
  o_2 <= slice1_y_net;
  o_3 <= slice2_y_net;
  o_4 <= slice3_y_net;
  o_5 <= slice4_y_net;
  o_6 <= slice5_y_net;
  o_7 <= slice6_y_net;
  o_8 <= slice7_y_net;
  o_9 <= slice8_y_net;
  o_10 <= slice9_y_net;
  o_11 <= slice10_y_net;
  o_12 <= slice11_y_net;
  o_13 <= slice12_y_net;
  o_14 <= slice13_y_net;
  o_15 <= slice14_y_net;
  o_16 <= slice15_y_net;
  bitbasher5_a_net <= i;
  slice0 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 15,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher5_a_net,
    y => slice0_y_net
  );
  slice1 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 16,
    new_msb => 31,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher5_a_net,
    y => slice1_y_net
  );
  slice2 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 32,
    new_msb => 47,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher5_a_net,
    y => slice2_y_net
  );
  slice3 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 48,
    new_msb => 63,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher5_a_net,
    y => slice3_y_net
  );
  slice4 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 64,
    new_msb => 79,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher5_a_net,
    y => slice4_y_net
  );
  slice5 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 80,
    new_msb => 95,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher5_a_net,
    y => slice5_y_net
  );
  slice6 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 96,
    new_msb => 111,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher5_a_net,
    y => slice6_y_net
  );
  slice7 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 112,
    new_msb => 127,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher5_a_net,
    y => slice7_y_net
  );
  slice8 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 128,
    new_msb => 143,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher5_a_net,
    y => slice8_y_net
  );
  slice9 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 144,
    new_msb => 159,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher5_a_net,
    y => slice9_y_net
  );
  slice10 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 160,
    new_msb => 175,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher5_a_net,
    y => slice10_y_net
  );
  slice11 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 176,
    new_msb => 191,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher5_a_net,
    y => slice11_y_net
  );
  slice12 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 192,
    new_msb => 207,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher5_a_net,
    y => slice12_y_net
  );
  slice13 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 208,
    new_msb => 223,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher5_a_net,
    y => slice13_y_net
  );
  slice14 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 224,
    new_msb => 239,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher5_a_net,
    y => slice14_y_net
  );
  slice15 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 240,
    new_msb => 255,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher5_a_net,
    y => slice15_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Scalar to Vector6
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_scalar_to_vector6 is
  port (
    i : in std_logic_vector( 256-1 downto 0 );
    o_1 : out std_logic_vector( 16-1 downto 0 );
    o_2 : out std_logic_vector( 16-1 downto 0 );
    o_3 : out std_logic_vector( 16-1 downto 0 );
    o_4 : out std_logic_vector( 16-1 downto 0 );
    o_5 : out std_logic_vector( 16-1 downto 0 );
    o_6 : out std_logic_vector( 16-1 downto 0 );
    o_7 : out std_logic_vector( 16-1 downto 0 );
    o_8 : out std_logic_vector( 16-1 downto 0 );
    o_9 : out std_logic_vector( 16-1 downto 0 );
    o_10 : out std_logic_vector( 16-1 downto 0 );
    o_11 : out std_logic_vector( 16-1 downto 0 );
    o_12 : out std_logic_vector( 16-1 downto 0 );
    o_13 : out std_logic_vector( 16-1 downto 0 );
    o_14 : out std_logic_vector( 16-1 downto 0 );
    o_15 : out std_logic_vector( 16-1 downto 0 );
    o_16 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_scalar_to_vector6;
architecture structural of psb3_0_scalar_to_vector6 is 
  signal slice7_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 16-1 downto 0 );
  signal bitbasher6_a_net : std_logic_vector( 256-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 16-1 downto 0 );
begin
  o_1 <= slice0_y_net;
  o_2 <= slice1_y_net;
  o_3 <= slice2_y_net;
  o_4 <= slice3_y_net;
  o_5 <= slice4_y_net;
  o_6 <= slice5_y_net;
  o_7 <= slice6_y_net;
  o_8 <= slice7_y_net;
  o_9 <= slice8_y_net;
  o_10 <= slice9_y_net;
  o_11 <= slice10_y_net;
  o_12 <= slice11_y_net;
  o_13 <= slice12_y_net;
  o_14 <= slice13_y_net;
  o_15 <= slice14_y_net;
  o_16 <= slice15_y_net;
  bitbasher6_a_net <= i;
  slice0 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 15,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher6_a_net,
    y => slice0_y_net
  );
  slice1 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 16,
    new_msb => 31,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher6_a_net,
    y => slice1_y_net
  );
  slice2 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 32,
    new_msb => 47,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher6_a_net,
    y => slice2_y_net
  );
  slice3 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 48,
    new_msb => 63,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher6_a_net,
    y => slice3_y_net
  );
  slice4 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 64,
    new_msb => 79,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher6_a_net,
    y => slice4_y_net
  );
  slice5 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 80,
    new_msb => 95,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher6_a_net,
    y => slice5_y_net
  );
  slice6 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 96,
    new_msb => 111,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher6_a_net,
    y => slice6_y_net
  );
  slice7 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 112,
    new_msb => 127,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher6_a_net,
    y => slice7_y_net
  );
  slice8 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 128,
    new_msb => 143,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher6_a_net,
    y => slice8_y_net
  );
  slice9 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 144,
    new_msb => 159,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher6_a_net,
    y => slice9_y_net
  );
  slice10 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 160,
    new_msb => 175,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher6_a_net,
    y => slice10_y_net
  );
  slice11 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 176,
    new_msb => 191,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher6_a_net,
    y => slice11_y_net
  );
  slice12 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 192,
    new_msb => 207,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher6_a_net,
    y => slice12_y_net
  );
  slice13 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 208,
    new_msb => 223,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher6_a_net,
    y => slice13_y_net
  );
  slice14 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 224,
    new_msb => 239,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher6_a_net,
    y => slice14_y_net
  );
  slice15 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 240,
    new_msb => 255,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher6_a_net,
    y => slice15_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Scalar to Vector7
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_scalar_to_vector7 is
  port (
    i : in std_logic_vector( 256-1 downto 0 );
    o_1 : out std_logic_vector( 16-1 downto 0 );
    o_2 : out std_logic_vector( 16-1 downto 0 );
    o_3 : out std_logic_vector( 16-1 downto 0 );
    o_4 : out std_logic_vector( 16-1 downto 0 );
    o_5 : out std_logic_vector( 16-1 downto 0 );
    o_6 : out std_logic_vector( 16-1 downto 0 );
    o_7 : out std_logic_vector( 16-1 downto 0 );
    o_8 : out std_logic_vector( 16-1 downto 0 );
    o_9 : out std_logic_vector( 16-1 downto 0 );
    o_10 : out std_logic_vector( 16-1 downto 0 );
    o_11 : out std_logic_vector( 16-1 downto 0 );
    o_12 : out std_logic_vector( 16-1 downto 0 );
    o_13 : out std_logic_vector( 16-1 downto 0 );
    o_14 : out std_logic_vector( 16-1 downto 0 );
    o_15 : out std_logic_vector( 16-1 downto 0 );
    o_16 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_scalar_to_vector7;
architecture structural of psb3_0_scalar_to_vector7 is 
  signal slice15_y_net : std_logic_vector( 16-1 downto 0 );
  signal bitbasher7_a_net : std_logic_vector( 256-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 16-1 downto 0 );
begin
  o_1 <= slice0_y_net;
  o_2 <= slice1_y_net;
  o_3 <= slice2_y_net;
  o_4 <= slice3_y_net;
  o_5 <= slice4_y_net;
  o_6 <= slice5_y_net;
  o_7 <= slice6_y_net;
  o_8 <= slice7_y_net;
  o_9 <= slice8_y_net;
  o_10 <= slice9_y_net;
  o_11 <= slice10_y_net;
  o_12 <= slice11_y_net;
  o_13 <= slice12_y_net;
  o_14 <= slice13_y_net;
  o_15 <= slice14_y_net;
  o_16 <= slice15_y_net;
  bitbasher7_a_net <= i;
  slice0 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 15,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher7_a_net,
    y => slice0_y_net
  );
  slice1 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 16,
    new_msb => 31,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher7_a_net,
    y => slice1_y_net
  );
  slice2 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 32,
    new_msb => 47,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher7_a_net,
    y => slice2_y_net
  );
  slice3 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 48,
    new_msb => 63,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher7_a_net,
    y => slice3_y_net
  );
  slice4 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 64,
    new_msb => 79,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher7_a_net,
    y => slice4_y_net
  );
  slice5 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 80,
    new_msb => 95,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher7_a_net,
    y => slice5_y_net
  );
  slice6 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 96,
    new_msb => 111,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher7_a_net,
    y => slice6_y_net
  );
  slice7 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 112,
    new_msb => 127,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher7_a_net,
    y => slice7_y_net
  );
  slice8 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 128,
    new_msb => 143,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher7_a_net,
    y => slice8_y_net
  );
  slice9 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 144,
    new_msb => 159,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher7_a_net,
    y => slice9_y_net
  );
  slice10 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 160,
    new_msb => 175,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher7_a_net,
    y => slice10_y_net
  );
  slice11 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 176,
    new_msb => 191,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher7_a_net,
    y => slice11_y_net
  );
  slice12 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 192,
    new_msb => 207,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher7_a_net,
    y => slice12_y_net
  );
  slice13 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 208,
    new_msb => 223,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher7_a_net,
    y => slice13_y_net
  );
  slice14 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 224,
    new_msb => 239,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher7_a_net,
    y => slice14_y_net
  );
  slice15 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 240,
    new_msb => 255,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher7_a_net,
    y => slice15_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Scalar to Vector8
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_scalar_to_vector8 is
  port (
    i : in std_logic_vector( 256-1 downto 0 );
    o_1 : out std_logic_vector( 16-1 downto 0 );
    o_2 : out std_logic_vector( 16-1 downto 0 );
    o_3 : out std_logic_vector( 16-1 downto 0 );
    o_4 : out std_logic_vector( 16-1 downto 0 );
    o_5 : out std_logic_vector( 16-1 downto 0 );
    o_6 : out std_logic_vector( 16-1 downto 0 );
    o_7 : out std_logic_vector( 16-1 downto 0 );
    o_8 : out std_logic_vector( 16-1 downto 0 );
    o_9 : out std_logic_vector( 16-1 downto 0 );
    o_10 : out std_logic_vector( 16-1 downto 0 );
    o_11 : out std_logic_vector( 16-1 downto 0 );
    o_12 : out std_logic_vector( 16-1 downto 0 );
    o_13 : out std_logic_vector( 16-1 downto 0 );
    o_14 : out std_logic_vector( 16-1 downto 0 );
    o_15 : out std_logic_vector( 16-1 downto 0 );
    o_16 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_scalar_to_vector8;
architecture structural of psb3_0_scalar_to_vector8 is 
  signal slice15_y_net : std_logic_vector( 16-1 downto 0 );
  signal bitbasher8_a_net : std_logic_vector( 256-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 16-1 downto 0 );
begin
  o_1 <= slice0_y_net;
  o_2 <= slice1_y_net;
  o_3 <= slice2_y_net;
  o_4 <= slice3_y_net;
  o_5 <= slice4_y_net;
  o_6 <= slice5_y_net;
  o_7 <= slice6_y_net;
  o_8 <= slice7_y_net;
  o_9 <= slice8_y_net;
  o_10 <= slice9_y_net;
  o_11 <= slice10_y_net;
  o_12 <= slice11_y_net;
  o_13 <= slice12_y_net;
  o_14 <= slice13_y_net;
  o_15 <= slice14_y_net;
  o_16 <= slice15_y_net;
  bitbasher8_a_net <= i;
  slice0 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 15,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher8_a_net,
    y => slice0_y_net
  );
  slice1 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 16,
    new_msb => 31,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher8_a_net,
    y => slice1_y_net
  );
  slice2 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 32,
    new_msb => 47,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher8_a_net,
    y => slice2_y_net
  );
  slice3 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 48,
    new_msb => 63,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher8_a_net,
    y => slice3_y_net
  );
  slice4 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 64,
    new_msb => 79,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher8_a_net,
    y => slice4_y_net
  );
  slice5 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 80,
    new_msb => 95,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher8_a_net,
    y => slice5_y_net
  );
  slice6 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 96,
    new_msb => 111,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher8_a_net,
    y => slice6_y_net
  );
  slice7 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 112,
    new_msb => 127,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher8_a_net,
    y => slice7_y_net
  );
  slice8 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 128,
    new_msb => 143,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher8_a_net,
    y => slice8_y_net
  );
  slice9 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 144,
    new_msb => 159,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher8_a_net,
    y => slice9_y_net
  );
  slice10 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 160,
    new_msb => 175,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher8_a_net,
    y => slice10_y_net
  );
  slice11 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 176,
    new_msb => 191,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher8_a_net,
    y => slice11_y_net
  );
  slice12 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 192,
    new_msb => 207,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher8_a_net,
    y => slice12_y_net
  );
  slice13 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 208,
    new_msb => 223,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher8_a_net,
    y => slice13_y_net
  );
  slice14 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 224,
    new_msb => 239,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher8_a_net,
    y => slice14_y_net
  );
  slice15 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 240,
    new_msb => 255,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => bitbasher8_a_net,
    y => slice15_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/ToneSelect/FIFO_delay
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_fifo_delay is
  port (
    in1 : in std_logic_vector( 16-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    out1 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_fifo_delay;
architecture structural of psb3_0_fifo_delay is 
  signal delay49_q_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret32_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal fifo3_full_net : std_logic;
  signal clk_net : std_logic;
  signal ce_net : std_logic;
  signal fifo3_empty_net : std_logic;
  signal constant17_op_net : std_logic_vector( 1-1 downto 0 );
  signal fifo3_dout_net : std_logic_vector( 16-1 downto 0 );
begin
  out1 <= fifo3_dout_net;
  reinterpret32_output_port_net <= in1;
  clk_net <= clk_1;
  ce_net <= ce_1;
  constant17 : entity xil_defaultlib.sysgen_constant_71e89d757c 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant17_op_net
  );
  delay49 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 261,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => constant17_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay49_q_net
  );
  fifo3 : entity xil_defaultlib.psb3_0_xlfifogen_u 
  generic map (
    core_name0 => "psb3_0_fifo_generator_i1",
    data_count_width => 10,
    data_width => 16,
    extra_registers => 1,
    has_ae => 0,
    has_af => 0,
    has_rst => false,
    ignore_din_for_gcd => false,
    percent_full_width => 1
  )
  port map (
    en => '1',
    rst => '0',
    din => reinterpret32_output_port_net,
    we => constant17_op_net(0),
    re => delay49_q_net(0),
    clk => clk_net,
    ce => ce_net,
    we_ce => ce_net,
    re_ce => ce_net,
    dout => fifo3_dout_net,
    empty => fifo3_empty_net,
    full => fifo3_full_net
  );
end structural;
-- Generated from Simulink block PSB3_0/ToneSelect/FIFO_delay1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_fifo_delay1 is
  port (
    in1 : in std_logic_vector( 16-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    out1 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_fifo_delay1;
architecture structural of psb3_0_fifo_delay1 is 
  signal reinterpret33_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal clk_net : std_logic;
  signal fifo3_dout_net : std_logic_vector( 16-1 downto 0 );
  signal ce_net : std_logic;
  signal fifo3_full_net : std_logic;
  signal constant17_op_net : std_logic_vector( 1-1 downto 0 );
  signal fifo3_empty_net : std_logic;
  signal delay49_q_net : std_logic_vector( 1-1 downto 0 );
begin
  out1 <= fifo3_dout_net;
  reinterpret33_output_port_net <= in1;
  clk_net <= clk_1;
  ce_net <= ce_1;
  constant17 : entity xil_defaultlib.sysgen_constant_71e89d757c 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant17_op_net
  );
  delay49 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 261,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => constant17_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay49_q_net
  );
  fifo3 : entity xil_defaultlib.psb3_0_xlfifogen_u 
  generic map (
    core_name0 => "psb3_0_fifo_generator_i1",
    data_count_width => 10,
    data_width => 16,
    extra_registers => 1,
    has_ae => 0,
    has_af => 0,
    has_rst => false,
    ignore_din_for_gcd => false,
    percent_full_width => 1
  )
  port map (
    en => '1',
    rst => '0',
    din => reinterpret33_output_port_net,
    we => constant17_op_net(0),
    re => delay49_q_net(0),
    clk => clk_net,
    ce => ce_net,
    we_ce => ce_net,
    re_ce => ce_net,
    dout => fifo3_dout_net,
    empty => fifo3_empty_net,
    full => fifo3_full_net
  );
end structural;
-- Generated from Simulink block PSB3_0/ToneSelect/FIFO_delay10
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_fifo_delay10 is
  port (
    in1 : in std_logic_vector( 16-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    out1 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_fifo_delay10;
architecture structural of psb3_0_fifo_delay10 is 
  signal fifo3_empty_net : std_logic;
  signal fifo3_full_net : std_logic;
  signal ce_net : std_logic;
  signal fifo3_dout_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret42_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal constant17_op_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal delay49_q_net : std_logic_vector( 1-1 downto 0 );
begin
  out1 <= fifo3_dout_net;
  reinterpret42_output_port_net <= in1;
  clk_net <= clk_1;
  ce_net <= ce_1;
  constant17 : entity xil_defaultlib.sysgen_constant_71e89d757c 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant17_op_net
  );
  delay49 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 261,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => constant17_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay49_q_net
  );
  fifo3 : entity xil_defaultlib.psb3_0_xlfifogen_u 
  generic map (
    core_name0 => "psb3_0_fifo_generator_i1",
    data_count_width => 10,
    data_width => 16,
    extra_registers => 1,
    has_ae => 0,
    has_af => 0,
    has_rst => false,
    ignore_din_for_gcd => false,
    percent_full_width => 1
  )
  port map (
    en => '1',
    rst => '0',
    din => reinterpret42_output_port_net,
    we => constant17_op_net(0),
    re => delay49_q_net(0),
    clk => clk_net,
    ce => ce_net,
    we_ce => ce_net,
    re_ce => ce_net,
    dout => fifo3_dout_net,
    empty => fifo3_empty_net,
    full => fifo3_full_net
  );
end structural;
-- Generated from Simulink block PSB3_0/ToneSelect/FIFO_delay11
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_fifo_delay11 is
  port (
    in1 : in std_logic_vector( 16-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    out1 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_fifo_delay11;
architecture structural of psb3_0_fifo_delay11 is 
  signal fifo3_dout_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret43_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal fifo3_full_net : std_logic;
  signal clk_net : std_logic;
  signal ce_net : std_logic;
  signal fifo3_empty_net : std_logic;
  signal delay49_q_net : std_logic_vector( 1-1 downto 0 );
  signal constant17_op_net : std_logic_vector( 1-1 downto 0 );
begin
  out1 <= fifo3_dout_net;
  reinterpret43_output_port_net <= in1;
  clk_net <= clk_1;
  ce_net <= ce_1;
  constant17 : entity xil_defaultlib.sysgen_constant_71e89d757c 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant17_op_net
  );
  delay49 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 261,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => constant17_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay49_q_net
  );
  fifo3 : entity xil_defaultlib.psb3_0_xlfifogen_u 
  generic map (
    core_name0 => "psb3_0_fifo_generator_i1",
    data_count_width => 10,
    data_width => 16,
    extra_registers => 1,
    has_ae => 0,
    has_af => 0,
    has_rst => false,
    ignore_din_for_gcd => false,
    percent_full_width => 1
  )
  port map (
    en => '1',
    rst => '0',
    din => reinterpret43_output_port_net,
    we => constant17_op_net(0),
    re => delay49_q_net(0),
    clk => clk_net,
    ce => ce_net,
    we_ce => ce_net,
    re_ce => ce_net,
    dout => fifo3_dout_net,
    empty => fifo3_empty_net,
    full => fifo3_full_net
  );
end structural;
-- Generated from Simulink block PSB3_0/ToneSelect/FIFO_delay12
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_fifo_delay12 is
  port (
    in1 : in std_logic_vector( 16-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    out1 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_fifo_delay12;
architecture structural of psb3_0_fifo_delay12 is 
  signal clk_net : std_logic;
  signal fifo3_dout_net : std_logic_vector( 16-1 downto 0 );
  signal constant17_op_net : std_logic_vector( 1-1 downto 0 );
  signal delay49_q_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret44_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal ce_net : std_logic;
  signal fifo3_empty_net : std_logic;
  signal fifo3_full_net : std_logic;
begin
  out1 <= fifo3_dout_net;
  reinterpret44_output_port_net <= in1;
  clk_net <= clk_1;
  ce_net <= ce_1;
  constant17 : entity xil_defaultlib.sysgen_constant_71e89d757c 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant17_op_net
  );
  delay49 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 261,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => constant17_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay49_q_net
  );
  fifo3 : entity xil_defaultlib.psb3_0_xlfifogen_u 
  generic map (
    core_name0 => "psb3_0_fifo_generator_i1",
    data_count_width => 10,
    data_width => 16,
    extra_registers => 1,
    has_ae => 0,
    has_af => 0,
    has_rst => false,
    ignore_din_for_gcd => false,
    percent_full_width => 1
  )
  port map (
    en => '1',
    rst => '0',
    din => reinterpret44_output_port_net,
    we => constant17_op_net(0),
    re => delay49_q_net(0),
    clk => clk_net,
    ce => ce_net,
    we_ce => ce_net,
    re_ce => ce_net,
    dout => fifo3_dout_net,
    empty => fifo3_empty_net,
    full => fifo3_full_net
  );
end structural;
-- Generated from Simulink block PSB3_0/ToneSelect/FIFO_delay13
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_fifo_delay13 is
  port (
    in1 : in std_logic_vector( 16-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    out1 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_fifo_delay13;
architecture structural of psb3_0_fifo_delay13 is 
  signal clk_net : std_logic;
  signal fifo3_full_net : std_logic;
  signal reinterpret45_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal ce_net : std_logic;
  signal delay49_q_net : std_logic_vector( 1-1 downto 0 );
  signal constant17_op_net : std_logic_vector( 1-1 downto 0 );
  signal fifo3_dout_net : std_logic_vector( 16-1 downto 0 );
  signal fifo3_empty_net : std_logic;
begin
  out1 <= fifo3_dout_net;
  reinterpret45_output_port_net <= in1;
  clk_net <= clk_1;
  ce_net <= ce_1;
  constant17 : entity xil_defaultlib.sysgen_constant_71e89d757c 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant17_op_net
  );
  delay49 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 261,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => constant17_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay49_q_net
  );
  fifo3 : entity xil_defaultlib.psb3_0_xlfifogen_u 
  generic map (
    core_name0 => "psb3_0_fifo_generator_i1",
    data_count_width => 10,
    data_width => 16,
    extra_registers => 1,
    has_ae => 0,
    has_af => 0,
    has_rst => false,
    ignore_din_for_gcd => false,
    percent_full_width => 1
  )
  port map (
    en => '1',
    rst => '0',
    din => reinterpret45_output_port_net,
    we => constant17_op_net(0),
    re => delay49_q_net(0),
    clk => clk_net,
    ce => ce_net,
    we_ce => ce_net,
    re_ce => ce_net,
    dout => fifo3_dout_net,
    empty => fifo3_empty_net,
    full => fifo3_full_net
  );
end structural;
-- Generated from Simulink block PSB3_0/ToneSelect/FIFO_delay14
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_fifo_delay14 is
  port (
    in1 : in std_logic_vector( 16-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    out1 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_fifo_delay14;
architecture structural of psb3_0_fifo_delay14 is 
  signal clk_net : std_logic;
  signal fifo3_dout_net : std_logic_vector( 16-1 downto 0 );
  signal constant17_op_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret46_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal delay49_q_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal fifo3_full_net : std_logic;
  signal fifo3_empty_net : std_logic;
begin
  out1 <= fifo3_dout_net;
  reinterpret46_output_port_net <= in1;
  clk_net <= clk_1;
  ce_net <= ce_1;
  constant17 : entity xil_defaultlib.sysgen_constant_71e89d757c 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant17_op_net
  );
  delay49 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 261,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => constant17_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay49_q_net
  );
  fifo3 : entity xil_defaultlib.psb3_0_xlfifogen_u 
  generic map (
    core_name0 => "psb3_0_fifo_generator_i1",
    data_count_width => 10,
    data_width => 16,
    extra_registers => 1,
    has_ae => 0,
    has_af => 0,
    has_rst => false,
    ignore_din_for_gcd => false,
    percent_full_width => 1
  )
  port map (
    en => '1',
    rst => '0',
    din => reinterpret46_output_port_net,
    we => constant17_op_net(0),
    re => delay49_q_net(0),
    clk => clk_net,
    ce => ce_net,
    we_ce => ce_net,
    re_ce => ce_net,
    dout => fifo3_dout_net,
    empty => fifo3_empty_net,
    full => fifo3_full_net
  );
end structural;
-- Generated from Simulink block PSB3_0/ToneSelect/FIFO_delay15
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_fifo_delay15 is
  port (
    in1 : in std_logic_vector( 16-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    out1 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_fifo_delay15;
architecture structural of psb3_0_fifo_delay15 is 
  signal fifo3_full_net : std_logic;
  signal clk_net : std_logic;
  signal ce_net : std_logic;
  signal fifo3_empty_net : std_logic;
  signal fifo3_dout_net : std_logic_vector( 16-1 downto 0 );
  signal delay49_q_net : std_logic_vector( 1-1 downto 0 );
  signal constant17_op_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret47_output_port_net : std_logic_vector( 16-1 downto 0 );
begin
  out1 <= fifo3_dout_net;
  reinterpret47_output_port_net <= in1;
  clk_net <= clk_1;
  ce_net <= ce_1;
  constant17 : entity xil_defaultlib.sysgen_constant_71e89d757c 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant17_op_net
  );
  delay49 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 261,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => constant17_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay49_q_net
  );
  fifo3 : entity xil_defaultlib.psb3_0_xlfifogen_u 
  generic map (
    core_name0 => "psb3_0_fifo_generator_i1",
    data_count_width => 10,
    data_width => 16,
    extra_registers => 1,
    has_ae => 0,
    has_af => 0,
    has_rst => false,
    ignore_din_for_gcd => false,
    percent_full_width => 1
  )
  port map (
    en => '1',
    rst => '0',
    din => reinterpret47_output_port_net,
    we => constant17_op_net(0),
    re => delay49_q_net(0),
    clk => clk_net,
    ce => ce_net,
    we_ce => ce_net,
    re_ce => ce_net,
    dout => fifo3_dout_net,
    empty => fifo3_empty_net,
    full => fifo3_full_net
  );
end structural;
-- Generated from Simulink block PSB3_0/ToneSelect/FIFO_delay2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_fifo_delay2 is
  port (
    in1 : in std_logic_vector( 16-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    out1 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_fifo_delay2;
architecture structural of psb3_0_fifo_delay2 is 
  signal fifo3_dout_net : std_logic_vector( 16-1 downto 0 );
  signal clk_net : std_logic;
  signal ce_net : std_logic;
  signal constant17_op_net : std_logic_vector( 1-1 downto 0 );
  signal delay49_q_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret34_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal fifo3_empty_net : std_logic;
  signal fifo3_full_net : std_logic;
begin
  out1 <= fifo3_dout_net;
  reinterpret34_output_port_net <= in1;
  clk_net <= clk_1;
  ce_net <= ce_1;
  constant17 : entity xil_defaultlib.sysgen_constant_71e89d757c 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant17_op_net
  );
  delay49 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 261,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => constant17_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay49_q_net
  );
  fifo3 : entity xil_defaultlib.psb3_0_xlfifogen_u 
  generic map (
    core_name0 => "psb3_0_fifo_generator_i1",
    data_count_width => 10,
    data_width => 16,
    extra_registers => 1,
    has_ae => 0,
    has_af => 0,
    has_rst => false,
    ignore_din_for_gcd => false,
    percent_full_width => 1
  )
  port map (
    en => '1',
    rst => '0',
    din => reinterpret34_output_port_net,
    we => constant17_op_net(0),
    re => delay49_q_net(0),
    clk => clk_net,
    ce => ce_net,
    we_ce => ce_net,
    re_ce => ce_net,
    dout => fifo3_dout_net,
    empty => fifo3_empty_net,
    full => fifo3_full_net
  );
end structural;
-- Generated from Simulink block PSB3_0/ToneSelect/FIFO_delay3
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_fifo_delay3 is
  port (
    in1 : in std_logic_vector( 16-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    out1 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_fifo_delay3;
architecture structural of psb3_0_fifo_delay3 is 
  signal ce_net : std_logic;
  signal reinterpret35_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal fifo3_empty_net : std_logic;
  signal fifo3_full_net : std_logic;
  signal delay49_q_net : std_logic_vector( 1-1 downto 0 );
  signal fifo3_dout_net : std_logic_vector( 16-1 downto 0 );
  signal clk_net : std_logic;
  signal constant17_op_net : std_logic_vector( 1-1 downto 0 );
begin
  out1 <= fifo3_dout_net;
  reinterpret35_output_port_net <= in1;
  clk_net <= clk_1;
  ce_net <= ce_1;
  constant17 : entity xil_defaultlib.sysgen_constant_71e89d757c 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant17_op_net
  );
  delay49 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 261,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => constant17_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay49_q_net
  );
  fifo3 : entity xil_defaultlib.psb3_0_xlfifogen_u 
  generic map (
    core_name0 => "psb3_0_fifo_generator_i1",
    data_count_width => 10,
    data_width => 16,
    extra_registers => 1,
    has_ae => 0,
    has_af => 0,
    has_rst => false,
    ignore_din_for_gcd => false,
    percent_full_width => 1
  )
  port map (
    en => '1',
    rst => '0',
    din => reinterpret35_output_port_net,
    we => constant17_op_net(0),
    re => delay49_q_net(0),
    clk => clk_net,
    ce => ce_net,
    we_ce => ce_net,
    re_ce => ce_net,
    dout => fifo3_dout_net,
    empty => fifo3_empty_net,
    full => fifo3_full_net
  );
end structural;
-- Generated from Simulink block PSB3_0/ToneSelect/FIFO_delay4
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_fifo_delay4 is
  port (
    in1 : in std_logic_vector( 16-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    out1 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_fifo_delay4;
architecture structural of psb3_0_fifo_delay4 is 
  signal reinterpret36_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal clk_net : std_logic;
  signal ce_net : std_logic;
  signal fifo3_dout_net : std_logic_vector( 16-1 downto 0 );
  signal constant17_op_net : std_logic_vector( 1-1 downto 0 );
  signal fifo3_full_net : std_logic;
  signal fifo3_empty_net : std_logic;
  signal delay49_q_net : std_logic_vector( 1-1 downto 0 );
begin
  out1 <= fifo3_dout_net;
  reinterpret36_output_port_net <= in1;
  clk_net <= clk_1;
  ce_net <= ce_1;
  constant17 : entity xil_defaultlib.sysgen_constant_71e89d757c 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant17_op_net
  );
  delay49 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 261,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => constant17_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay49_q_net
  );
  fifo3 : entity xil_defaultlib.psb3_0_xlfifogen_u 
  generic map (
    core_name0 => "psb3_0_fifo_generator_i1",
    data_count_width => 10,
    data_width => 16,
    extra_registers => 1,
    has_ae => 0,
    has_af => 0,
    has_rst => false,
    ignore_din_for_gcd => false,
    percent_full_width => 1
  )
  port map (
    en => '1',
    rst => '0',
    din => reinterpret36_output_port_net,
    we => constant17_op_net(0),
    re => delay49_q_net(0),
    clk => clk_net,
    ce => ce_net,
    we_ce => ce_net,
    re_ce => ce_net,
    dout => fifo3_dout_net,
    empty => fifo3_empty_net,
    full => fifo3_full_net
  );
end structural;
-- Generated from Simulink block PSB3_0/ToneSelect/FIFO_delay5
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_fifo_delay5 is
  port (
    in1 : in std_logic_vector( 16-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    out1 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_fifo_delay5;
architecture structural of psb3_0_fifo_delay5 is 
  signal ce_net : std_logic;
  signal fifo3_empty_net : std_logic;
  signal fifo3_full_net : std_logic;
  signal reinterpret37_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal fifo3_dout_net : std_logic_vector( 16-1 downto 0 );
  signal delay49_q_net : std_logic_vector( 1-1 downto 0 );
  signal constant17_op_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
begin
  out1 <= fifo3_dout_net;
  reinterpret37_output_port_net <= in1;
  clk_net <= clk_1;
  ce_net <= ce_1;
  constant17 : entity xil_defaultlib.sysgen_constant_71e89d757c 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant17_op_net
  );
  delay49 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 261,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => constant17_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay49_q_net
  );
  fifo3 : entity xil_defaultlib.psb3_0_xlfifogen_u 
  generic map (
    core_name0 => "psb3_0_fifo_generator_i1",
    data_count_width => 10,
    data_width => 16,
    extra_registers => 1,
    has_ae => 0,
    has_af => 0,
    has_rst => false,
    ignore_din_for_gcd => false,
    percent_full_width => 1
  )
  port map (
    en => '1',
    rst => '0',
    din => reinterpret37_output_port_net,
    we => constant17_op_net(0),
    re => delay49_q_net(0),
    clk => clk_net,
    ce => ce_net,
    we_ce => ce_net,
    re_ce => ce_net,
    dout => fifo3_dout_net,
    empty => fifo3_empty_net,
    full => fifo3_full_net
  );
end structural;
-- Generated from Simulink block PSB3_0/ToneSelect/FIFO_delay6
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_fifo_delay6 is
  port (
    in1 : in std_logic_vector( 16-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    out1 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_fifo_delay6;
architecture structural of psb3_0_fifo_delay6 is 
  signal fifo3_dout_net : std_logic_vector( 16-1 downto 0 );
  signal clk_net : std_logic;
  signal ce_net : std_logic;
  signal reinterpret38_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal fifo3_empty_net : std_logic;
  signal constant17_op_net : std_logic_vector( 1-1 downto 0 );
  signal delay49_q_net : std_logic_vector( 1-1 downto 0 );
  signal fifo3_full_net : std_logic;
begin
  out1 <= fifo3_dout_net;
  reinterpret38_output_port_net <= in1;
  clk_net <= clk_1;
  ce_net <= ce_1;
  constant17 : entity xil_defaultlib.sysgen_constant_71e89d757c 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant17_op_net
  );
  delay49 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 261,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => constant17_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay49_q_net
  );
  fifo3 : entity xil_defaultlib.psb3_0_xlfifogen_u 
  generic map (
    core_name0 => "psb3_0_fifo_generator_i1",
    data_count_width => 10,
    data_width => 16,
    extra_registers => 1,
    has_ae => 0,
    has_af => 0,
    has_rst => false,
    ignore_din_for_gcd => false,
    percent_full_width => 1
  )
  port map (
    en => '1',
    rst => '0',
    din => reinterpret38_output_port_net,
    we => constant17_op_net(0),
    re => delay49_q_net(0),
    clk => clk_net,
    ce => ce_net,
    we_ce => ce_net,
    re_ce => ce_net,
    dout => fifo3_dout_net,
    empty => fifo3_empty_net,
    full => fifo3_full_net
  );
end structural;
-- Generated from Simulink block PSB3_0/ToneSelect/FIFO_delay7
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_fifo_delay7 is
  port (
    in1 : in std_logic_vector( 16-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    out1 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_fifo_delay7;
architecture structural of psb3_0_fifo_delay7 is 
  signal fifo3_full_net : std_logic;
  signal fifo3_empty_net : std_logic;
  signal constant17_op_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret39_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal clk_net : std_logic;
  signal delay49_q_net : std_logic_vector( 1-1 downto 0 );
  signal fifo3_dout_net : std_logic_vector( 16-1 downto 0 );
  signal ce_net : std_logic;
begin
  out1 <= fifo3_dout_net;
  reinterpret39_output_port_net <= in1;
  clk_net <= clk_1;
  ce_net <= ce_1;
  constant17 : entity xil_defaultlib.sysgen_constant_71e89d757c 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant17_op_net
  );
  delay49 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 261,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => constant17_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay49_q_net
  );
  fifo3 : entity xil_defaultlib.psb3_0_xlfifogen_u 
  generic map (
    core_name0 => "psb3_0_fifo_generator_i1",
    data_count_width => 10,
    data_width => 16,
    extra_registers => 1,
    has_ae => 0,
    has_af => 0,
    has_rst => false,
    ignore_din_for_gcd => false,
    percent_full_width => 1
  )
  port map (
    en => '1',
    rst => '0',
    din => reinterpret39_output_port_net,
    we => constant17_op_net(0),
    re => delay49_q_net(0),
    clk => clk_net,
    ce => ce_net,
    we_ce => ce_net,
    re_ce => ce_net,
    dout => fifo3_dout_net,
    empty => fifo3_empty_net,
    full => fifo3_full_net
  );
end structural;
-- Generated from Simulink block PSB3_0/ToneSelect/FIFO_delay8
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_fifo_delay8 is
  port (
    in1 : in std_logic_vector( 16-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    out1 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_fifo_delay8;
architecture structural of psb3_0_fifo_delay8 is 
  signal fifo3_full_net : std_logic;
  signal fifo3_dout_net : std_logic_vector( 16-1 downto 0 );
  signal clk_net : std_logic;
  signal ce_net : std_logic;
  signal delay49_q_net : std_logic_vector( 1-1 downto 0 );
  signal constant17_op_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret40_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal fifo3_empty_net : std_logic;
begin
  out1 <= fifo3_dout_net;
  reinterpret40_output_port_net <= in1;
  clk_net <= clk_1;
  ce_net <= ce_1;
  constant17 : entity xil_defaultlib.sysgen_constant_71e89d757c 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant17_op_net
  );
  delay49 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 261,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => constant17_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay49_q_net
  );
  fifo3 : entity xil_defaultlib.psb3_0_xlfifogen_u 
  generic map (
    core_name0 => "psb3_0_fifo_generator_i1",
    data_count_width => 10,
    data_width => 16,
    extra_registers => 1,
    has_ae => 0,
    has_af => 0,
    has_rst => false,
    ignore_din_for_gcd => false,
    percent_full_width => 1
  )
  port map (
    en => '1',
    rst => '0',
    din => reinterpret40_output_port_net,
    we => constant17_op_net(0),
    re => delay49_q_net(0),
    clk => clk_net,
    ce => ce_net,
    we_ce => ce_net,
    re_ce => ce_net,
    dout => fifo3_dout_net,
    empty => fifo3_empty_net,
    full => fifo3_full_net
  );
end structural;
-- Generated from Simulink block PSB3_0/ToneSelect/FIFO_delay9
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_fifo_delay9 is
  port (
    in1 : in std_logic_vector( 16-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    out1 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_fifo_delay9;
architecture structural of psb3_0_fifo_delay9 is 
  signal clk_net : std_logic;
  signal reinterpret41_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal ce_net : std_logic;
  signal constant17_op_net : std_logic_vector( 1-1 downto 0 );
  signal fifo3_dout_net : std_logic_vector( 16-1 downto 0 );
  signal fifo3_full_net : std_logic;
  signal delay49_q_net : std_logic_vector( 1-1 downto 0 );
  signal fifo3_empty_net : std_logic;
begin
  out1 <= fifo3_dout_net;
  reinterpret41_output_port_net <= in1;
  clk_net <= clk_1;
  ce_net <= ce_1;
  constant17 : entity xil_defaultlib.sysgen_constant_71e89d757c 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant17_op_net
  );
  delay49 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 261,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => constant17_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay49_q_net
  );
  fifo3 : entity xil_defaultlib.psb3_0_xlfifogen_u 
  generic map (
    core_name0 => "psb3_0_fifo_generator_i1",
    data_count_width => 10,
    data_width => 16,
    extra_registers => 1,
    has_ae => 0,
    has_af => 0,
    has_rst => false,
    ignore_din_for_gcd => false,
    percent_full_width => 1
  )
  port map (
    en => '1',
    rst => '0',
    din => reinterpret41_output_port_net,
    we => constant17_op_net(0),
    re => delay49_q_net(0),
    clk => clk_net,
    ce => ce_net,
    we_ce => ce_net,
    re_ce => ce_net,
    dout => fifo3_dout_net,
    empty => fifo3_empty_net,
    full => fifo3_full_net
  );
end structural;
-- Generated from Simulink block PSB3_0/ToneSelect/imag_slice_0
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_imag_slice_0 is
  port (
    sel : in std_logic_vector( 3-1 downto 0 );
    input : in std_logic_vector( 256-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    output : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_imag_slice_0;
architecture structural of psb3_0_imag_slice_0 is 
  signal mux1_y_net : std_logic_vector( 256-1 downto 0 );
  signal mux20_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 16-1 downto 0 );
  signal clk_net : std_logic;
  signal slice8_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 16-1 downto 0 );
  signal ce_net : std_logic;
  signal parallel_sel_0_y_net : std_logic_vector( 3-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 16-1 downto 0 );
begin
  output <= mux20_y_net;
  parallel_sel_0_y_net <= sel;
  mux1_y_net <= input;
  clk_net <= clk_1;
  ce_net <= ce_1;
  mux20 : entity xil_defaultlib.sysgen_mux_f12f18e758 
  port map (
    clr => '0',
    sel => parallel_sel_0_y_net,
    d0 => slice2_y_net,
    d1 => slice1_y_net,
    d2 => slice3_y_net,
    d3 => slice4_y_net,
    d4 => slice5_y_net,
    d5 => slice6_y_net,
    d6 => slice7_y_net,
    d7 => slice8_y_net,
    clk => clk_net,
    ce => ce_net,
    y => mux20_y_net
  );
  slice1 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 48,
    new_msb => 63,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux1_y_net,
    y => slice1_y_net
  );
  slice2 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 16,
    new_msb => 31,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux1_y_net,
    y => slice2_y_net
  );
  slice3 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 80,
    new_msb => 95,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux1_y_net,
    y => slice3_y_net
  );
  slice4 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 112,
    new_msb => 127,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux1_y_net,
    y => slice4_y_net
  );
  slice5 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 144,
    new_msb => 159,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux1_y_net,
    y => slice5_y_net
  );
  slice6 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 176,
    new_msb => 191,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux1_y_net,
    y => slice6_y_net
  );
  slice7 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 208,
    new_msb => 223,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux1_y_net,
    y => slice7_y_net
  );
  slice8 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 240,
    new_msb => 255,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux1_y_net,
    y => slice8_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/ToneSelect/imag_slice_1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_imag_slice_1 is
  port (
    sel : in std_logic_vector( 3-1 downto 0 );
    input : in std_logic_vector( 256-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    output : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_imag_slice_1;
architecture structural of psb3_0_imag_slice_1 is 
  signal slice6_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 16-1 downto 0 );
  signal ce_net : std_logic;
  signal mux20_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 16-1 downto 0 );
  signal mux20_y_net_x0 : std_logic_vector( 256-1 downto 0 );
  signal clk_net : std_logic;
  signal slice5_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 16-1 downto 0 );
  signal parallel_sel_1_y_net : std_logic_vector( 3-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 16-1 downto 0 );
begin
  output <= mux20_y_net;
  parallel_sel_1_y_net <= sel;
  mux20_y_net_x0 <= input;
  clk_net <= clk_1;
  ce_net <= ce_1;
  mux20 : entity xil_defaultlib.sysgen_mux_f12f18e758 
  port map (
    clr => '0',
    sel => parallel_sel_1_y_net,
    d0 => slice2_y_net,
    d1 => slice1_y_net,
    d2 => slice3_y_net,
    d3 => slice4_y_net,
    d4 => slice5_y_net,
    d5 => slice6_y_net,
    d6 => slice7_y_net,
    d7 => slice8_y_net,
    clk => clk_net,
    ce => ce_net,
    y => mux20_y_net
  );
  slice1 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 48,
    new_msb => 63,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux20_y_net_x0,
    y => slice1_y_net
  );
  slice2 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 16,
    new_msb => 31,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux20_y_net_x0,
    y => slice2_y_net
  );
  slice3 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 80,
    new_msb => 95,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux20_y_net_x0,
    y => slice3_y_net
  );
  slice4 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 112,
    new_msb => 127,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux20_y_net_x0,
    y => slice4_y_net
  );
  slice5 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 144,
    new_msb => 159,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux20_y_net_x0,
    y => slice5_y_net
  );
  slice6 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 176,
    new_msb => 191,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux20_y_net_x0,
    y => slice6_y_net
  );
  slice7 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 208,
    new_msb => 223,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux20_y_net_x0,
    y => slice7_y_net
  );
  slice8 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 240,
    new_msb => 255,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux20_y_net_x0,
    y => slice8_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/ToneSelect/imag_slice_2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_imag_slice_2 is
  port (
    sel : in std_logic_vector( 3-1 downto 0 );
    input : in std_logic_vector( 256-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    output : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_imag_slice_2;
architecture structural of psb3_0_imag_slice_2 is 
  signal mux20_y_net : std_logic_vector( 16-1 downto 0 );
  signal ce_net : std_logic;
  signal mux21_y_net : std_logic_vector( 256-1 downto 0 );
  signal clk_net : std_logic;
  signal parallel_sel_2_y_net : std_logic_vector( 3-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 16-1 downto 0 );
begin
  output <= mux20_y_net;
  parallel_sel_2_y_net <= sel;
  mux21_y_net <= input;
  clk_net <= clk_1;
  ce_net <= ce_1;
  mux20 : entity xil_defaultlib.sysgen_mux_f12f18e758 
  port map (
    clr => '0',
    sel => parallel_sel_2_y_net,
    d0 => slice2_y_net,
    d1 => slice1_y_net,
    d2 => slice3_y_net,
    d3 => slice4_y_net,
    d4 => slice5_y_net,
    d5 => slice6_y_net,
    d6 => slice7_y_net,
    d7 => slice8_y_net,
    clk => clk_net,
    ce => ce_net,
    y => mux20_y_net
  );
  slice1 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 48,
    new_msb => 63,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux21_y_net,
    y => slice1_y_net
  );
  slice2 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 16,
    new_msb => 31,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux21_y_net,
    y => slice2_y_net
  );
  slice3 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 80,
    new_msb => 95,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux21_y_net,
    y => slice3_y_net
  );
  slice4 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 112,
    new_msb => 127,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux21_y_net,
    y => slice4_y_net
  );
  slice5 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 144,
    new_msb => 159,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux21_y_net,
    y => slice5_y_net
  );
  slice6 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 176,
    new_msb => 191,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux21_y_net,
    y => slice6_y_net
  );
  slice7 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 208,
    new_msb => 223,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux21_y_net,
    y => slice7_y_net
  );
  slice8 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 240,
    new_msb => 255,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux21_y_net,
    y => slice8_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/ToneSelect/imag_slice_3
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_imag_slice_3 is
  port (
    sel : in std_logic_vector( 3-1 downto 0 );
    input : in std_logic_vector( 256-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    output : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_imag_slice_3;
architecture structural of psb3_0_imag_slice_3 is 
  signal slice4_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 16-1 downto 0 );
  signal ce_net : std_logic;
  signal mux20_y_net : std_logic_vector( 16-1 downto 0 );
  signal clk_net : std_logic;
  signal parallel_sel_3_y_net : std_logic_vector( 3-1 downto 0 );
  signal mux22_y_net : std_logic_vector( 256-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 16-1 downto 0 );
begin
  output <= mux20_y_net;
  parallel_sel_3_y_net <= sel;
  mux22_y_net <= input;
  clk_net <= clk_1;
  ce_net <= ce_1;
  mux20 : entity xil_defaultlib.sysgen_mux_f12f18e758 
  port map (
    clr => '0',
    sel => parallel_sel_3_y_net,
    d0 => slice2_y_net,
    d1 => slice1_y_net,
    d2 => slice3_y_net,
    d3 => slice4_y_net,
    d4 => slice5_y_net,
    d5 => slice6_y_net,
    d6 => slice7_y_net,
    d7 => slice8_y_net,
    clk => clk_net,
    ce => ce_net,
    y => mux20_y_net
  );
  slice1 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 48,
    new_msb => 63,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux22_y_net,
    y => slice1_y_net
  );
  slice2 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 16,
    new_msb => 31,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux22_y_net,
    y => slice2_y_net
  );
  slice3 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 80,
    new_msb => 95,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux22_y_net,
    y => slice3_y_net
  );
  slice4 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 112,
    new_msb => 127,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux22_y_net,
    y => slice4_y_net
  );
  slice5 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 144,
    new_msb => 159,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux22_y_net,
    y => slice5_y_net
  );
  slice6 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 176,
    new_msb => 191,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux22_y_net,
    y => slice6_y_net
  );
  slice7 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 208,
    new_msb => 223,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux22_y_net,
    y => slice7_y_net
  );
  slice8 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 240,
    new_msb => 255,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux22_y_net,
    y => slice8_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/ToneSelect/imag_slice_4
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_imag_slice_4 is
  port (
    sel : in std_logic_vector( 3-1 downto 0 );
    input : in std_logic_vector( 256-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    output : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_imag_slice_4;
architecture structural of psb3_0_imag_slice_4 is 
  signal parallel_sel_4_y_net : std_logic_vector( 3-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 16-1 downto 0 );
  signal clk_net : std_logic;
  signal slice5_y_net : std_logic_vector( 16-1 downto 0 );
  signal ce_net : std_logic;
  signal slice1_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 16-1 downto 0 );
  signal mux23_y_net : std_logic_vector( 256-1 downto 0 );
  signal mux20_y_net : std_logic_vector( 16-1 downto 0 );
begin
  output <= mux20_y_net;
  parallel_sel_4_y_net <= sel;
  mux23_y_net <= input;
  clk_net <= clk_1;
  ce_net <= ce_1;
  mux20 : entity xil_defaultlib.sysgen_mux_f12f18e758 
  port map (
    clr => '0',
    sel => parallel_sel_4_y_net,
    d0 => slice2_y_net,
    d1 => slice1_y_net,
    d2 => slice3_y_net,
    d3 => slice4_y_net,
    d4 => slice5_y_net,
    d5 => slice6_y_net,
    d6 => slice7_y_net,
    d7 => slice8_y_net,
    clk => clk_net,
    ce => ce_net,
    y => mux20_y_net
  );
  slice1 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 48,
    new_msb => 63,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux23_y_net,
    y => slice1_y_net
  );
  slice2 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 16,
    new_msb => 31,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux23_y_net,
    y => slice2_y_net
  );
  slice3 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 80,
    new_msb => 95,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux23_y_net,
    y => slice3_y_net
  );
  slice4 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 112,
    new_msb => 127,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux23_y_net,
    y => slice4_y_net
  );
  slice5 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 144,
    new_msb => 159,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux23_y_net,
    y => slice5_y_net
  );
  slice6 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 176,
    new_msb => 191,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux23_y_net,
    y => slice6_y_net
  );
  slice7 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 208,
    new_msb => 223,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux23_y_net,
    y => slice7_y_net
  );
  slice8 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 240,
    new_msb => 255,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux23_y_net,
    y => slice8_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/ToneSelect/imag_slice_5
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_imag_slice_5 is
  port (
    sel : in std_logic_vector( 3-1 downto 0 );
    input : in std_logic_vector( 256-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    output : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_imag_slice_5;
architecture structural of psb3_0_imag_slice_5 is 
  signal slice1_y_net : std_logic_vector( 16-1 downto 0 );
  signal ce_net : std_logic;
  signal slice3_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 16-1 downto 0 );
  signal parallel_sel_5_y_net : std_logic_vector( 3-1 downto 0 );
  signal mux24_y_net : std_logic_vector( 256-1 downto 0 );
  signal clk_net : std_logic;
  signal slice8_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 16-1 downto 0 );
  signal mux20_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 16-1 downto 0 );
begin
  output <= mux20_y_net;
  parallel_sel_5_y_net <= sel;
  mux24_y_net <= input;
  clk_net <= clk_1;
  ce_net <= ce_1;
  mux20 : entity xil_defaultlib.sysgen_mux_f12f18e758 
  port map (
    clr => '0',
    sel => parallel_sel_5_y_net,
    d0 => slice2_y_net,
    d1 => slice1_y_net,
    d2 => slice3_y_net,
    d3 => slice4_y_net,
    d4 => slice5_y_net,
    d5 => slice6_y_net,
    d6 => slice7_y_net,
    d7 => slice8_y_net,
    clk => clk_net,
    ce => ce_net,
    y => mux20_y_net
  );
  slice1 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 48,
    new_msb => 63,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux24_y_net,
    y => slice1_y_net
  );
  slice2 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 16,
    new_msb => 31,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux24_y_net,
    y => slice2_y_net
  );
  slice3 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 80,
    new_msb => 95,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux24_y_net,
    y => slice3_y_net
  );
  slice4 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 112,
    new_msb => 127,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux24_y_net,
    y => slice4_y_net
  );
  slice5 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 144,
    new_msb => 159,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux24_y_net,
    y => slice5_y_net
  );
  slice6 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 176,
    new_msb => 191,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux24_y_net,
    y => slice6_y_net
  );
  slice7 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 208,
    new_msb => 223,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux24_y_net,
    y => slice7_y_net
  );
  slice8 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 240,
    new_msb => 255,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux24_y_net,
    y => slice8_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/ToneSelect/imag_slice_6
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_imag_slice_6 is
  port (
    sel : in std_logic_vector( 3-1 downto 0 );
    input : in std_logic_vector( 256-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    output : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_imag_slice_6;
architecture structural of psb3_0_imag_slice_6 is 
  signal mux25_y_net : std_logic_vector( 256-1 downto 0 );
  signal mux20_y_net : std_logic_vector( 16-1 downto 0 );
  signal clk_net : std_logic;
  signal parallel_sel_6_y_net : std_logic_vector( 3-1 downto 0 );
  signal ce_net : std_logic;
  signal slice5_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 16-1 downto 0 );
begin
  output <= mux20_y_net;
  parallel_sel_6_y_net <= sel;
  mux25_y_net <= input;
  clk_net <= clk_1;
  ce_net <= ce_1;
  mux20 : entity xil_defaultlib.sysgen_mux_f12f18e758 
  port map (
    clr => '0',
    sel => parallel_sel_6_y_net,
    d0 => slice2_y_net,
    d1 => slice1_y_net,
    d2 => slice3_y_net,
    d3 => slice4_y_net,
    d4 => slice5_y_net,
    d5 => slice6_y_net,
    d6 => slice7_y_net,
    d7 => slice8_y_net,
    clk => clk_net,
    ce => ce_net,
    y => mux20_y_net
  );
  slice1 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 48,
    new_msb => 63,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux25_y_net,
    y => slice1_y_net
  );
  slice2 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 16,
    new_msb => 31,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux25_y_net,
    y => slice2_y_net
  );
  slice3 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 80,
    new_msb => 95,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux25_y_net,
    y => slice3_y_net
  );
  slice4 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 112,
    new_msb => 127,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux25_y_net,
    y => slice4_y_net
  );
  slice5 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 144,
    new_msb => 159,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux25_y_net,
    y => slice5_y_net
  );
  slice6 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 176,
    new_msb => 191,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux25_y_net,
    y => slice6_y_net
  );
  slice7 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 208,
    new_msb => 223,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux25_y_net,
    y => slice7_y_net
  );
  slice8 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 240,
    new_msb => 255,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux25_y_net,
    y => slice8_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/ToneSelect/imag_slice_7
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_imag_slice_7 is
  port (
    sel : in std_logic_vector( 3-1 downto 0 );
    input : in std_logic_vector( 256-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    output : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_imag_slice_7;
architecture structural of psb3_0_imag_slice_7 is 
  signal parallel_sel_7_y_net : std_logic_vector( 3-1 downto 0 );
  signal mux20_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 16-1 downto 0 );
  signal ce_net : std_logic;
  signal clk_net : std_logic;
  signal slice2_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 16-1 downto 0 );
  signal mux26_y_net : std_logic_vector( 256-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 16-1 downto 0 );
begin
  output <= mux20_y_net;
  parallel_sel_7_y_net <= sel;
  mux26_y_net <= input;
  clk_net <= clk_1;
  ce_net <= ce_1;
  mux20 : entity xil_defaultlib.sysgen_mux_f12f18e758 
  port map (
    clr => '0',
    sel => parallel_sel_7_y_net,
    d0 => slice2_y_net,
    d1 => slice1_y_net,
    d2 => slice3_y_net,
    d3 => slice4_y_net,
    d4 => slice5_y_net,
    d5 => slice6_y_net,
    d6 => slice7_y_net,
    d7 => slice8_y_net,
    clk => clk_net,
    ce => ce_net,
    y => mux20_y_net
  );
  slice1 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 48,
    new_msb => 63,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux26_y_net,
    y => slice1_y_net
  );
  slice2 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 16,
    new_msb => 31,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux26_y_net,
    y => slice2_y_net
  );
  slice3 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 80,
    new_msb => 95,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux26_y_net,
    y => slice3_y_net
  );
  slice4 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 112,
    new_msb => 127,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux26_y_net,
    y => slice4_y_net
  );
  slice5 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 144,
    new_msb => 159,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux26_y_net,
    y => slice5_y_net
  );
  slice6 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 176,
    new_msb => 191,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux26_y_net,
    y => slice6_y_net
  );
  slice7 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 208,
    new_msb => 223,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux26_y_net,
    y => slice7_y_net
  );
  slice8 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 240,
    new_msb => 255,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux26_y_net,
    y => slice8_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/ToneSelect/real_slice_0
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_real_slice_0 is
  port (
    sel : in std_logic_vector( 3-1 downto 0 );
    input : in std_logic_vector( 256-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    output : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_real_slice_0;
architecture structural of psb3_0_real_slice_0 is 
  signal mux1_y_net : std_logic_vector( 256-1 downto 0 );
  signal mux20_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 16-1 downto 0 );
  signal parallel_sel_0_y_net : std_logic_vector( 3-1 downto 0 );
  signal clk_net : std_logic;
  signal slice4_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 16-1 downto 0 );
  signal ce_net : std_logic;
begin
  output <= mux20_y_net;
  parallel_sel_0_y_net <= sel;
  mux1_y_net <= input;
  clk_net <= clk_1;
  ce_net <= ce_1;
  mux20 : entity xil_defaultlib.sysgen_mux_f12f18e758 
  port map (
    clr => '0',
    sel => parallel_sel_0_y_net,
    d0 => slice2_y_net,
    d1 => slice1_y_net,
    d2 => slice3_y_net,
    d3 => slice4_y_net,
    d4 => slice5_y_net,
    d5 => slice6_y_net,
    d6 => slice7_y_net,
    d7 => slice8_y_net,
    clk => clk_net,
    ce => ce_net,
    y => mux20_y_net
  );
  slice1 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 32,
    new_msb => 47,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux1_y_net,
    y => slice1_y_net
  );
  slice2 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 15,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux1_y_net,
    y => slice2_y_net
  );
  slice3 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 64,
    new_msb => 79,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux1_y_net,
    y => slice3_y_net
  );
  slice4 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 96,
    new_msb => 111,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux1_y_net,
    y => slice4_y_net
  );
  slice5 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 128,
    new_msb => 143,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux1_y_net,
    y => slice5_y_net
  );
  slice6 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 160,
    new_msb => 175,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux1_y_net,
    y => slice6_y_net
  );
  slice7 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 192,
    new_msb => 207,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux1_y_net,
    y => slice7_y_net
  );
  slice8 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 224,
    new_msb => 239,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux1_y_net,
    y => slice8_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/ToneSelect/real_slice_1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_real_slice_1 is
  port (
    sel : in std_logic_vector( 3-1 downto 0 );
    input : in std_logic_vector( 256-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    output : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_real_slice_1;
architecture structural of psb3_0_real_slice_1 is 
  signal slice6_y_net : std_logic_vector( 16-1 downto 0 );
  signal clk_net : std_logic;
  signal slice5_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 16-1 downto 0 );
  signal mux20_y_net : std_logic_vector( 16-1 downto 0 );
  signal parallel_sel_1_y_net : std_logic_vector( 3-1 downto 0 );
  signal mux20_y_net_x0 : std_logic_vector( 256-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 16-1 downto 0 );
  signal ce_net : std_logic;
  signal slice2_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 16-1 downto 0 );
begin
  output <= mux20_y_net;
  parallel_sel_1_y_net <= sel;
  mux20_y_net_x0 <= input;
  clk_net <= clk_1;
  ce_net <= ce_1;
  mux20 : entity xil_defaultlib.sysgen_mux_f12f18e758 
  port map (
    clr => '0',
    sel => parallel_sel_1_y_net,
    d0 => slice2_y_net,
    d1 => slice1_y_net,
    d2 => slice3_y_net,
    d3 => slice4_y_net,
    d4 => slice5_y_net,
    d5 => slice6_y_net,
    d6 => slice7_y_net,
    d7 => slice8_y_net,
    clk => clk_net,
    ce => ce_net,
    y => mux20_y_net
  );
  slice1 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 32,
    new_msb => 47,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux20_y_net_x0,
    y => slice1_y_net
  );
  slice2 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 15,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux20_y_net_x0,
    y => slice2_y_net
  );
  slice3 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 64,
    new_msb => 79,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux20_y_net_x0,
    y => slice3_y_net
  );
  slice4 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 96,
    new_msb => 111,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux20_y_net_x0,
    y => slice4_y_net
  );
  slice5 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 128,
    new_msb => 143,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux20_y_net_x0,
    y => slice5_y_net
  );
  slice6 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 160,
    new_msb => 175,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux20_y_net_x0,
    y => slice6_y_net
  );
  slice7 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 192,
    new_msb => 207,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux20_y_net_x0,
    y => slice7_y_net
  );
  slice8 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 224,
    new_msb => 239,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux20_y_net_x0,
    y => slice8_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/ToneSelect/real_slice_2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_real_slice_2 is
  port (
    sel : in std_logic_vector( 3-1 downto 0 );
    input : in std_logic_vector( 256-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    output : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_real_slice_2;
architecture structural of psb3_0_real_slice_2 is 
  signal mux20_y_net : std_logic_vector( 16-1 downto 0 );
  signal parallel_sel_2_y_net : std_logic_vector( 3-1 downto 0 );
  signal mux21_y_net : std_logic_vector( 256-1 downto 0 );
  signal clk_net : std_logic;
  signal ce_net : std_logic;
  signal slice1_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 16-1 downto 0 );
begin
  output <= mux20_y_net;
  parallel_sel_2_y_net <= sel;
  mux21_y_net <= input;
  clk_net <= clk_1;
  ce_net <= ce_1;
  mux20 : entity xil_defaultlib.sysgen_mux_f12f18e758 
  port map (
    clr => '0',
    sel => parallel_sel_2_y_net,
    d0 => slice2_y_net,
    d1 => slice1_y_net,
    d2 => slice3_y_net,
    d3 => slice4_y_net,
    d4 => slice5_y_net,
    d5 => slice6_y_net,
    d6 => slice7_y_net,
    d7 => slice8_y_net,
    clk => clk_net,
    ce => ce_net,
    y => mux20_y_net
  );
  slice1 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 32,
    new_msb => 47,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux21_y_net,
    y => slice1_y_net
  );
  slice2 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 15,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux21_y_net,
    y => slice2_y_net
  );
  slice3 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 64,
    new_msb => 79,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux21_y_net,
    y => slice3_y_net
  );
  slice4 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 96,
    new_msb => 111,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux21_y_net,
    y => slice4_y_net
  );
  slice5 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 128,
    new_msb => 143,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux21_y_net,
    y => slice5_y_net
  );
  slice6 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 160,
    new_msb => 175,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux21_y_net,
    y => slice6_y_net
  );
  slice7 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 192,
    new_msb => 207,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux21_y_net,
    y => slice7_y_net
  );
  slice8 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 224,
    new_msb => 239,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux21_y_net,
    y => slice8_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/ToneSelect/real_slice_3
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_real_slice_3 is
  port (
    sel : in std_logic_vector( 3-1 downto 0 );
    input : in std_logic_vector( 256-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    output : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_real_slice_3;
architecture structural of psb3_0_real_slice_3 is 
  signal parallel_sel_3_y_net : std_logic_vector( 3-1 downto 0 );
  signal mux20_y_net : std_logic_vector( 16-1 downto 0 );
  signal mux22_y_net : std_logic_vector( 256-1 downto 0 );
  signal ce_net : std_logic;
  signal clk_net : std_logic;
  signal slice2_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 16-1 downto 0 );
begin
  output <= mux20_y_net;
  parallel_sel_3_y_net <= sel;
  mux22_y_net <= input;
  clk_net <= clk_1;
  ce_net <= ce_1;
  mux20 : entity xil_defaultlib.sysgen_mux_f12f18e758 
  port map (
    clr => '0',
    sel => parallel_sel_3_y_net,
    d0 => slice2_y_net,
    d1 => slice1_y_net,
    d2 => slice3_y_net,
    d3 => slice4_y_net,
    d4 => slice5_y_net,
    d5 => slice6_y_net,
    d6 => slice7_y_net,
    d7 => slice8_y_net,
    clk => clk_net,
    ce => ce_net,
    y => mux20_y_net
  );
  slice1 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 32,
    new_msb => 47,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux22_y_net,
    y => slice1_y_net
  );
  slice2 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 15,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux22_y_net,
    y => slice2_y_net
  );
  slice3 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 64,
    new_msb => 79,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux22_y_net,
    y => slice3_y_net
  );
  slice4 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 96,
    new_msb => 111,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux22_y_net,
    y => slice4_y_net
  );
  slice5 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 128,
    new_msb => 143,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux22_y_net,
    y => slice5_y_net
  );
  slice6 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 160,
    new_msb => 175,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux22_y_net,
    y => slice6_y_net
  );
  slice7 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 192,
    new_msb => 207,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux22_y_net,
    y => slice7_y_net
  );
  slice8 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 224,
    new_msb => 239,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux22_y_net,
    y => slice8_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/ToneSelect/real_slice_4
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_real_slice_4 is
  port (
    sel : in std_logic_vector( 3-1 downto 0 );
    input : in std_logic_vector( 256-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    output : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_real_slice_4;
architecture structural of psb3_0_real_slice_4 is 
  signal mux23_y_net : std_logic_vector( 256-1 downto 0 );
  signal clk_net : std_logic;
  signal slice4_y_net : std_logic_vector( 16-1 downto 0 );
  signal ce_net : std_logic;
  signal slice7_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 16-1 downto 0 );
  signal mux20_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 16-1 downto 0 );
  signal parallel_sel_4_y_net : std_logic_vector( 3-1 downto 0 );
begin
  output <= mux20_y_net;
  parallel_sel_4_y_net <= sel;
  mux23_y_net <= input;
  clk_net <= clk_1;
  ce_net <= ce_1;
  mux20 : entity xil_defaultlib.sysgen_mux_f12f18e758 
  port map (
    clr => '0',
    sel => parallel_sel_4_y_net,
    d0 => slice2_y_net,
    d1 => slice1_y_net,
    d2 => slice3_y_net,
    d3 => slice4_y_net,
    d4 => slice5_y_net,
    d5 => slice6_y_net,
    d6 => slice7_y_net,
    d7 => slice8_y_net,
    clk => clk_net,
    ce => ce_net,
    y => mux20_y_net
  );
  slice1 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 32,
    new_msb => 47,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux23_y_net,
    y => slice1_y_net
  );
  slice2 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 15,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux23_y_net,
    y => slice2_y_net
  );
  slice3 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 64,
    new_msb => 79,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux23_y_net,
    y => slice3_y_net
  );
  slice4 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 96,
    new_msb => 111,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux23_y_net,
    y => slice4_y_net
  );
  slice5 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 128,
    new_msb => 143,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux23_y_net,
    y => slice5_y_net
  );
  slice6 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 160,
    new_msb => 175,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux23_y_net,
    y => slice6_y_net
  );
  slice7 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 192,
    new_msb => 207,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux23_y_net,
    y => slice7_y_net
  );
  slice8 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 224,
    new_msb => 239,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux23_y_net,
    y => slice8_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/ToneSelect/real_slice_5
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_real_slice_5 is
  port (
    sel : in std_logic_vector( 3-1 downto 0 );
    input : in std_logic_vector( 256-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    output : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_real_slice_5;
architecture structural of psb3_0_real_slice_5 is 
  signal clk_net : std_logic;
  signal slice2_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 16-1 downto 0 );
  signal mux24_y_net : std_logic_vector( 256-1 downto 0 );
  signal ce_net : std_logic;
  signal slice6_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 16-1 downto 0 );
  signal parallel_sel_5_y_net : std_logic_vector( 3-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 16-1 downto 0 );
  signal mux20_y_net : std_logic_vector( 16-1 downto 0 );
begin
  output <= mux20_y_net;
  parallel_sel_5_y_net <= sel;
  mux24_y_net <= input;
  clk_net <= clk_1;
  ce_net <= ce_1;
  mux20 : entity xil_defaultlib.sysgen_mux_f12f18e758 
  port map (
    clr => '0',
    sel => parallel_sel_5_y_net,
    d0 => slice2_y_net,
    d1 => slice1_y_net,
    d2 => slice3_y_net,
    d3 => slice4_y_net,
    d4 => slice5_y_net,
    d5 => slice6_y_net,
    d6 => slice7_y_net,
    d7 => slice8_y_net,
    clk => clk_net,
    ce => ce_net,
    y => mux20_y_net
  );
  slice1 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 32,
    new_msb => 47,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux24_y_net,
    y => slice1_y_net
  );
  slice2 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 15,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux24_y_net,
    y => slice2_y_net
  );
  slice3 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 64,
    new_msb => 79,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux24_y_net,
    y => slice3_y_net
  );
  slice4 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 96,
    new_msb => 111,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux24_y_net,
    y => slice4_y_net
  );
  slice5 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 128,
    new_msb => 143,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux24_y_net,
    y => slice5_y_net
  );
  slice6 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 160,
    new_msb => 175,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux24_y_net,
    y => slice6_y_net
  );
  slice7 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 192,
    new_msb => 207,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux24_y_net,
    y => slice7_y_net
  );
  slice8 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 224,
    new_msb => 239,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux24_y_net,
    y => slice8_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/ToneSelect/real_slice_6
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_real_slice_6 is
  port (
    sel : in std_logic_vector( 3-1 downto 0 );
    input : in std_logic_vector( 256-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    output : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_real_slice_6;
architecture structural of psb3_0_real_slice_6 is 
  signal mux20_y_net : std_logic_vector( 16-1 downto 0 );
  signal clk_net : std_logic;
  signal ce_net : std_logic;
  signal parallel_sel_6_y_net : std_logic_vector( 3-1 downto 0 );
  signal mux25_y_net : std_logic_vector( 256-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 16-1 downto 0 );
begin
  output <= mux20_y_net;
  parallel_sel_6_y_net <= sel;
  mux25_y_net <= input;
  clk_net <= clk_1;
  ce_net <= ce_1;
  mux20 : entity xil_defaultlib.sysgen_mux_f12f18e758 
  port map (
    clr => '0',
    sel => parallel_sel_6_y_net,
    d0 => slice2_y_net,
    d1 => slice1_y_net,
    d2 => slice3_y_net,
    d3 => slice4_y_net,
    d4 => slice5_y_net,
    d5 => slice6_y_net,
    d6 => slice7_y_net,
    d7 => slice8_y_net,
    clk => clk_net,
    ce => ce_net,
    y => mux20_y_net
  );
  slice1 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 32,
    new_msb => 47,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux25_y_net,
    y => slice1_y_net
  );
  slice2 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 15,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux25_y_net,
    y => slice2_y_net
  );
  slice3 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 64,
    new_msb => 79,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux25_y_net,
    y => slice3_y_net
  );
  slice4 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 96,
    new_msb => 111,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux25_y_net,
    y => slice4_y_net
  );
  slice5 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 128,
    new_msb => 143,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux25_y_net,
    y => slice5_y_net
  );
  slice6 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 160,
    new_msb => 175,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux25_y_net,
    y => slice6_y_net
  );
  slice7 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 192,
    new_msb => 207,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux25_y_net,
    y => slice7_y_net
  );
  slice8 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 224,
    new_msb => 239,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux25_y_net,
    y => slice8_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/ToneSelect/real_slice_7
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_real_slice_7 is
  port (
    sel : in std_logic_vector( 3-1 downto 0 );
    input : in std_logic_vector( 256-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    output : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_real_slice_7;
architecture structural of psb3_0_real_slice_7 is 
  signal mux26_y_net : std_logic_vector( 256-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 16-1 downto 0 );
  signal parallel_sel_7_y_net : std_logic_vector( 3-1 downto 0 );
  signal clk_net : std_logic;
  signal ce_net : std_logic;
  signal slice1_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 16-1 downto 0 );
  signal mux20_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 16-1 downto 0 );
begin
  output <= mux20_y_net;
  parallel_sel_7_y_net <= sel;
  mux26_y_net <= input;
  clk_net <= clk_1;
  ce_net <= ce_1;
  mux20 : entity xil_defaultlib.sysgen_mux_f12f18e758 
  port map (
    clr => '0',
    sel => parallel_sel_7_y_net,
    d0 => slice2_y_net,
    d1 => slice1_y_net,
    d2 => slice3_y_net,
    d3 => slice4_y_net,
    d4 => slice5_y_net,
    d5 => slice6_y_net,
    d6 => slice7_y_net,
    d7 => slice8_y_net,
    clk => clk_net,
    ce => ce_net,
    y => mux20_y_net
  );
  slice1 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 32,
    new_msb => 47,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux26_y_net,
    y => slice1_y_net
  );
  slice2 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 15,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux26_y_net,
    y => slice2_y_net
  );
  slice3 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 64,
    new_msb => 79,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux26_y_net,
    y => slice3_y_net
  );
  slice4 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 96,
    new_msb => 111,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux26_y_net,
    y => slice4_y_net
  );
  slice5 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 128,
    new_msb => 143,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux26_y_net,
    y => slice5_y_net
  );
  slice6 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 160,
    new_msb => 175,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux26_y_net,
    y => slice6_y_net
  );
  slice7 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 192,
    new_msb => 207,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux26_y_net,
    y => slice7_y_net
  );
  slice8 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 224,
    new_msb => 239,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux26_y_net,
    y => slice8_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/ToneSelect
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_toneselect is
  port (
    in_even1_im : in std_logic_vector( 16-1 downto 0 );
    in_even1_re : in std_logic_vector( 16-1 downto 0 );
    in_odd1_im : in std_logic_vector( 16-1 downto 0 );
    in_odd1_re : in std_logic_vector( 16-1 downto 0 );
    in_even2_im : in std_logic_vector( 16-1 downto 0 );
    in_even2_re : in std_logic_vector( 16-1 downto 0 );
    in_odd2_im : in std_logic_vector( 16-1 downto 0 );
    in_odd2_re : in std_logic_vector( 16-1 downto 0 );
    in_even3_im : in std_logic_vector( 16-1 downto 0 );
    in_even3_re : in std_logic_vector( 16-1 downto 0 );
    in_odd3_im : in std_logic_vector( 16-1 downto 0 );
    in_odd3_re : in std_logic_vector( 16-1 downto 0 );
    in_even4_im : in std_logic_vector( 16-1 downto 0 );
    in_even4_re : in std_logic_vector( 16-1 downto 0 );
    in_odd4_im : in std_logic_vector( 16-1 downto 0 );
    in_odd4_re : in std_logic_vector( 16-1 downto 0 );
    in_tvalid : in std_logic;
    rst : in std_logic_vector( 1-1 downto 0 );
    data_0 : in std_logic_vector( 12-1 downto 0 );
    data_1 : in std_logic_vector( 12-1 downto 0 );
    data_2 : in std_logic_vector( 12-1 downto 0 );
    data_3 : in std_logic_vector( 12-1 downto 0 );
    data_4 : in std_logic_vector( 12-1 downto 0 );
    data_5 : in std_logic_vector( 12-1 downto 0 );
    data_6 : in std_logic_vector( 12-1 downto 0 );
    data_7 : in std_logic_vector( 12-1 downto 0 );
    w_addr_x0 : in std_logic_vector( 8-1 downto 0 );
    we : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    out_even1_re : out std_logic_vector( 17-1 downto 0 );
    out_odd1_re : out std_logic_vector( 17-1 downto 0 );
    out_even2_re : out std_logic_vector( 17-1 downto 0 );
    out_odd2_re : out std_logic_vector( 17-1 downto 0 );
    out_even3_re : out std_logic_vector( 17-1 downto 0 );
    out_odd3_re : out std_logic_vector( 17-1 downto 0 );
    out_even4_re : out std_logic_vector( 17-1 downto 0 );
    out_odd4_re : out std_logic_vector( 17-1 downto 0 );
    out_even1_im : out std_logic_vector( 17-1 downto 0 );
    out_odd1_im : out std_logic_vector( 17-1 downto 0 );
    out_even2_im : out std_logic_vector( 17-1 downto 0 );
    out_odd2_im : out std_logic_vector( 17-1 downto 0 );
    out_even3_im : out std_logic_vector( 17-1 downto 0 );
    out_odd3_im : out std_logic_vector( 17-1 downto 0 );
    out_even4_im : out std_logic_vector( 17-1 downto 0 );
    out_odd4_im : out std_logic_vector( 17-1 downto 0 );
    out_tvalid : out std_logic_vector( 1-1 downto 0 )
  );
end psb3_0_toneselect;
architecture structural of psb3_0_toneselect is 
  signal bitbasher7_o_net : std_logic_vector( 17-1 downto 0 );
  signal bitbasher9_o_net : std_logic_vector( 17-1 downto 0 );
  signal bitbasher14_o_net : std_logic_vector( 17-1 downto 0 );
  signal bitbasher4_o_net : std_logic_vector( 17-1 downto 0 );
  signal bitbasher8_o_net : std_logic_vector( 17-1 downto 0 );
  signal bitbasher13_o_net : std_logic_vector( 17-1 downto 0 );
  signal bitbasher2_o_net : std_logic_vector( 17-1 downto 0 );
  signal bitbasher15_o_net : std_logic_vector( 17-1 downto 0 );
  signal bitbasher3_o_net : std_logic_vector( 17-1 downto 0 );
  signal bitbasher5_o_net : std_logic_vector( 17-1 downto 0 );
  signal bitbasher6_o_net : std_logic_vector( 17-1 downto 0 );
  signal constant14_op_net : std_logic_vector( 3-1 downto 0 );
  signal constant_op_net : std_logic_vector( 17-1 downto 0 );
  signal constant15_op_net : std_logic_vector( 17-1 downto 0 );
  signal constant16_op_net : std_logic_vector( 3-1 downto 0 );
  signal constant12_op_net : std_logic_vector( 3-1 downto 0 );
  signal constant10_op_net : std_logic_vector( 3-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 3-1 downto 0 );
  signal concat_y_net : std_logic_vector( 256-1 downto 0 );
  signal constant11_op_net : std_logic_vector( 17-1 downto 0 );
  signal constant13_op_net : std_logic_vector( 17-1 downto 0 );
  signal constant3_op_net : std_logic_vector( 17-1 downto 0 );
  signal constant7_op_net : std_logic_vector( 17-1 downto 0 );
  signal constant5_op_net : std_logic_vector( 17-1 downto 0 );
  signal convert_dout_net : std_logic_vector( 1-1 downto 0 );
  signal constant8_op_net : std_logic_vector( 3-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 12-1 downto 0 );
  signal constant4_op_net : std_logic_vector( 3-1 downto 0 );
  signal constant6_op_net : std_logic_vector( 3-1 downto 0 );
  signal constant9_op_net : std_logic_vector( 17-1 downto 0 );
  signal counter1_op_net : std_logic_vector( 8-1 downto 0 );
  signal constant2_op_net : std_logic_vector( 8-1 downto 0 );
  signal single_port_ram17_data_out_net : std_logic_vector( 12-1 downto 0 );
  signal mux29_y_net : std_logic_vector( 17-1 downto 0 );
  signal mux30_y_net : std_logic_vector( 17-1 downto 0 );
  signal mux2_y_net : std_logic_vector( 17-1 downto 0 );
  signal mux37_y_net : std_logic_vector( 17-1 downto 0 );
  signal mux33_y_net : std_logic_vector( 17-1 downto 0 );
  signal mux38_y_net : std_logic_vector( 17-1 downto 0 );
  signal mux42_y_net : std_logic_vector( 17-1 downto 0 );
  signal mux34_y_net : std_logic_vector( 17-1 downto 0 );
  signal mux46_y_net : std_logic_vector( 17-1 downto 0 );
  signal mux50_y_net : std_logic_vector( 17-1 downto 0 );
  signal delay11_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal cordic_6_0_even_1_m_axis_dout_tdata_imag_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal cordic_6_0_even_1_m_axis_dout_tdata_real_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal mux45_y_net : std_logic_vector( 17-1 downto 0 );
  signal mux54_y_net : std_logic_vector( 17-1 downto 0 );
  signal mux49_y_net : std_logic_vector( 17-1 downto 0 );
  signal cordic_6_0_odd_1_m_axis_dout_tdata_real_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal mux53_y_net : std_logic_vector( 17-1 downto 0 );
  signal cordic_6_0_odd_1_m_axis_dout_tdata_imag_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal cordic_6_0_even_2_m_axis_dout_tdata_imag_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal mux41_y_net : std_logic_vector( 17-1 downto 0 );
  signal cordic_6_0_even_2_m_axis_dout_tdata_real_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal mux27_y_net : std_logic_vector( 17-1 downto 0 );
  signal delay12_q_net : std_logic_vector( 8-1 downto 0 );
  signal fifo3_dout_net_x11 : std_logic_vector( 16-1 downto 0 );
  signal gin_tl_reset_net : std_logic_vector( 1-1 downto 0 );
  signal cordic_6_0_odd_2_m_axis_dout_tdata_real_net : std_logic_vector( 16-1 downto 0 );
  signal cordic_6_0_odd_1_m_axis_dout_tdata_imag_net : std_logic_vector( 16-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 12-1 downto 0 );
  signal cordic_6_0_even_1_m_axis_dout_tvalid_net : std_logic;
  signal delay9_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay7_q_net : std_logic_vector( 12-1 downto 0 );
  signal cordic_6_0_even_2_m_axis_dout_tdata_real_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret32_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret45_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret46_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal cordic_6_0_even_1_m_axis_dout_tdata_real_net : std_logic_vector( 16-1 downto 0 );
  signal fifo3_dout_net_x7 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret47_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal cordic_6_0_odd_1_m_axis_dout_tdata_real_net : std_logic_vector( 16-1 downto 0 );
  signal cordic_6_0_even_2_m_axis_dout_tdata_imag_net : std_logic_vector( 16-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 12-1 downto 0 );
  signal cordic_6_0_odd_2_m_axis_dout_tdata_imag_net : std_logic_vector( 16-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 12-1 downto 0 );
  signal ce_net : std_logic;
  signal delay11_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay16_q_net : std_logic_vector( 1-1 downto 0 );
  signal fifo3_dout_net_x13 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret33_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal fifo3_dout_net_x12 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret42_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret43_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal cordic_6_0_odd_2_m_axis_dout_tdata_real_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal fifo3_dout_net_x10 : std_logic_vector( 16-1 downto 0 );
  signal cordic_6_0_even_1_m_axis_dout_tdata_imag_net : std_logic_vector( 16-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay10_q_net : std_logic_vector( 12-1 downto 0 );
  signal reinterpret44_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal fifo3_dout_net_x8 : std_logic_vector( 16-1 downto 0 );
  signal clk_net : std_logic;
  signal fifo3_dout_net_x14 : std_logic_vector( 16-1 downto 0 );
  signal cordic_6_0_odd_2_m_axis_dout_tdata_imag_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal fifo3_dout_net_x9 : std_logic_vector( 16-1 downto 0 );
  signal parallel_sel_2_y_net : std_logic_vector( 3-1 downto 0 );
  signal fifo3_dout_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal parallel_sel_3_y_net : std_logic_vector( 3-1 downto 0 );
  signal mux20_y_net_x3 : std_logic_vector( 16-1 downto 0 );
  signal mux20_y_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal mux20_y_net_x13 : std_logic_vector( 16-1 downto 0 );
  signal mux22_y_net : std_logic_vector( 256-1 downto 0 );
  signal mux24_y_net : std_logic_vector( 256-1 downto 0 );
  signal parallel_sel_5_y_net : std_logic_vector( 3-1 downto 0 );
  signal reinterpret41_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal relational1_op_net : std_logic_vector( 1-1 downto 0 );
  signal mux20_y_net_x4 : std_logic_vector( 16-1 downto 0 );
  signal delay13_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 256-1 downto 0 );
  signal mux20_y_net_x1 : std_logic_vector( 16-1 downto 0 );
  signal mux26_y_net : std_logic_vector( 256-1 downto 0 );
  signal parallel_sel_0_y_net : std_logic_vector( 3-1 downto 0 );
  signal parallel_sel_6_y_net : std_logic_vector( 3-1 downto 0 );
  signal mux20_y_net_x14 : std_logic_vector( 16-1 downto 0 );
  signal fifo3_dout_net_x2 : std_logic_vector( 16-1 downto 0 );
  signal parallel_sel_7_y_net : std_logic_vector( 3-1 downto 0 );
  signal mux20_y_net_x2 : std_logic_vector( 16-1 downto 0 );
  signal fifo3_dout_net : std_logic_vector( 16-1 downto 0 );
  signal mux20_y_net_x7 : std_logic_vector( 16-1 downto 0 );
  signal accumulator_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux20_y_net_x6 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret34_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal fifo3_dout_net_x6 : std_logic_vector( 16-1 downto 0 );
  signal mux20_y_net_x8 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret35_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal fifo3_dout_net_x4 : std_logic_vector( 16-1 downto 0 );
  signal mux21_y_net : std_logic_vector( 256-1 downto 0 );
  signal reinterpret37_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mux20_y_net_x5 : std_logic_vector( 16-1 downto 0 );
  signal mux20_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret39_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal parallel_sel_4_y_net : std_logic_vector( 3-1 downto 0 );
  signal mux23_y_net : std_logic_vector( 256-1 downto 0 );
  signal mux20_y_net_x12 : std_logic_vector( 16-1 downto 0 );
  signal mux20_y_net_x10 : std_logic_vector( 16-1 downto 0 );
  signal mux20_y_net_x9 : std_logic_vector( 16-1 downto 0 );
  signal fifo3_dout_net_x5 : std_logic_vector( 16-1 downto 0 );
  signal mux25_y_net : std_logic_vector( 256-1 downto 0 );
  signal reinterpret38_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal parallel_sel_1_y_net : std_logic_vector( 3-1 downto 0 );
  signal mux20_y_net_x11 : std_logic_vector( 16-1 downto 0 );
  signal mux20_y_net_x15 : std_logic_vector( 256-1 downto 0 );
  signal reinterpret36_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal fifo3_dout_net_x3 : std_logic_vector( 16-1 downto 0 );
  signal fifo3_dout_net_x1 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret40_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub13_s_net : std_logic_vector( 17-1 downto 0 );
  signal reinterpret25_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret21_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret28_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub10_s_net : std_logic_vector( 17-1 downto 0 );
  signal reinterpret29_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret22_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 17-1 downto 0 );
  signal addsub11_s_net : std_logic_vector( 17-1 downto 0 );
  signal reinterpret23_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret24_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret27_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret20_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub12_s_net : std_logic_vector( 17-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub_s_net : std_logic_vector( 17-1 downto 0 );
  signal reinterpret26_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub14_s_net : std_logic_vector( 17-1 downto 0 );
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret31_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub5_s_net : std_logic_vector( 17-1 downto 0 );
  signal addsub15_s_net : std_logic_vector( 17-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub3_s_net : std_logic_vector( 17-1 downto 0 );
  signal addsub6_s_net : std_logic_vector( 17-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret30_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 17-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 17-1 downto 0 );
  signal reinterpret16_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub9_s_net : std_logic_vector( 17-1 downto 0 );
  signal reinterpret17_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal bitbasher_o_net : std_logic_vector( 17-1 downto 0 );
  signal addsub8_s_net : std_logic_vector( 17-1 downto 0 );
  signal bitbasher12_o_net : std_logic_vector( 17-1 downto 0 );
  signal bitbasher10_o_net : std_logic_vector( 17-1 downto 0 );
  signal addsub7_s_net : std_logic_vector( 17-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret19_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal bitbasher1_o_net : std_logic_vector( 17-1 downto 0 );
  signal reinterpret18_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal bitbasher11_o_net : std_logic_vector( 17-1 downto 0 );
  signal delay14_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay15_q_net : std_logic_vector( 8-1 downto 0 );
  signal delay12_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay17_q_net : std_logic_vector( 8-1 downto 0 );
  signal delay18_q_net : std_logic_vector( 1-1 downto 0 );
  signal bypass_bool_1_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay16_q_net_x0 : std_logic_vector( 8-1 downto 0 );
  signal addr_0_y_net : std_logic_vector( 8-1 downto 0 );
  signal bypass_bool_0_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay10_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal addr_2_y_net : std_logic_vector( 8-1 downto 0 );
  signal delay21_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay22_q_net : std_logic_vector( 8-1 downto 0 );
  signal delay25_q_net : std_logic_vector( 8-1 downto 0 );
  signal addr_1_y_net : std_logic_vector( 8-1 downto 0 );
  signal delay19_q_net : std_logic_vector( 8-1 downto 0 );
  signal delay20_q_net : std_logic_vector( 8-1 downto 0 );
  signal bypass_bool_2_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay23_q_net : std_logic_vector( 8-1 downto 0 );
  signal delay24_q_net : std_logic_vector( 1-1 downto 0 );
  signal bypass_bool_3_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net_x0 : std_logic_vector( 256-1 downto 0 );
  signal delay27_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay29_q_net : std_logic_vector( 8-1 downto 0 );
  signal addr_4_y_net : std_logic_vector( 8-1 downto 0 );
  signal single_port_ram18_data_out_net : std_logic_vector( 12-1 downto 0 );
  signal delay3_q_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal delay26_q_net : std_logic_vector( 8-1 downto 0 );
  signal delay31_q_net : std_logic_vector( 8-1 downto 0 );
  signal delay30_q_net : std_logic_vector( 1-1 downto 0 );
  signal bypass_bool_4_y_net : std_logic_vector( 1-1 downto 0 );
  signal addr_5_y_net : std_logic_vector( 8-1 downto 0 );
  signal delay32_q_net : std_logic_vector( 8-1 downto 0 );
  signal addr_3_y_net : std_logic_vector( 8-1 downto 0 );
  signal bypass_bool_5_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay28_q_net : std_logic_vector( 8-1 downto 0 );
  signal delay33_q_net : std_logic_vector( 1-1 downto 0 );
  signal bypass_bool_6_y_net : std_logic_vector( 1-1 downto 0 );
  signal single_port_ram19_data_out_net : std_logic_vector( 12-1 downto 0 );
  signal single_port_ram20_data_out_net : std_logic_vector( 12-1 downto 0 );
  signal addr_7_y_net : std_logic_vector( 8-1 downto 0 );
  signal delay5_q_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal delay38_q_net : std_logic_vector( 8-1 downto 0 );
  signal delay4_q_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal delay35_q_net : std_logic_vector( 8-1 downto 0 );
  signal addr_6_y_net : std_logic_vector( 8-1 downto 0 );
  signal delay36_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay37_q_net : std_logic_vector( 8-1 downto 0 );
  signal bypass_bool_7_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay39_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay34_q_net : std_logic_vector( 8-1 downto 0 );
  signal delay9_q_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal single_port_ram24_data_out_net : std_logic_vector( 12-1 downto 0 );
  signal inverter_op_net : std_logic_vector( 1-1 downto 0 );
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
  signal relational2_op_net : std_logic_vector( 1-1 downto 0 );
  signal relational_op_net : std_logic_vector( 1-1 downto 0 );
  signal logical1_y_net : std_logic_vector( 1-1 downto 0 );
  signal relational6_op_net : std_logic_vector( 1-1 downto 0 );
  signal single_port_ram22_data_out_net : std_logic_vector( 12-1 downto 0 );
  signal delay7_q_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal single_port_ram23_data_out_net : std_logic_vector( 12-1 downto 0 );
  signal relational3_op_net : std_logic_vector( 1-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 12-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 12-1 downto 0 );
  signal logical2_y_net : std_logic_vector( 1-1 downto 0 );
  signal relational4_op_net : std_logic_vector( 1-1 downto 0 );
  signal relational5_op_net : std_logic_vector( 1-1 downto 0 );
  signal single_port_ram21_data_out_net : std_logic_vector( 12-1 downto 0 );
  signal relational9_op_net : std_logic_vector( 1-1 downto 0 );
  signal relational8_op_net : std_logic_vector( 1-1 downto 0 );
  signal relational16_op_net : std_logic_vector( 1-1 downto 0 );
  signal logical5_y_net : std_logic_vector( 1-1 downto 0 );
  signal logical6_y_net : std_logic_vector( 1-1 downto 0 );
  signal relational11_op_net : std_logic_vector( 1-1 downto 0 );
  signal relational13_op_net : std_logic_vector( 1-1 downto 0 );
  signal relational10_op_net : std_logic_vector( 1-1 downto 0 );
  signal relational7_op_net : std_logic_vector( 1-1 downto 0 );
  signal logical4_y_net : std_logic_vector( 1-1 downto 0 );
  signal single_port_ram1_data_out_net : std_logic_vector( 256-1 downto 0 );
  signal logical3_y_net : std_logic_vector( 1-1 downto 0 );
  signal logical7_y_net : std_logic_vector( 1-1 downto 0 );
  signal relational15_op_net : std_logic_vector( 1-1 downto 0 );
  signal relational12_op_net : std_logic_vector( 1-1 downto 0 );
  signal relational14_op_net : std_logic_vector( 1-1 downto 0 );
  signal single_port_ram9_data_out_net : std_logic_vector( 256-1 downto 0 );
  signal mux10_y_net : std_logic_vector( 8-1 downto 0 );
  signal mux12_y_net : std_logic_vector( 8-1 downto 0 );
  signal mux11_y_net : std_logic_vector( 8-1 downto 0 );
  signal mux16_y_net : std_logic_vector( 8-1 downto 0 );
  signal mux17_y_net : std_logic_vector( 8-1 downto 0 );
  signal mux18_y_net : std_logic_vector( 8-1 downto 0 );
  signal mux13_y_net : std_logic_vector( 8-1 downto 0 );
  signal mux14_y_net : std_logic_vector( 8-1 downto 0 );
  signal mux15_y_net : std_logic_vector( 8-1 downto 0 );
  signal single_port_ram12_data_out_net : std_logic_vector( 256-1 downto 0 );
  signal single_port_ram2_data_out_net : std_logic_vector( 256-1 downto 0 );
  signal single_port_ram14_data_out_net : std_logic_vector( 256-1 downto 0 );
  signal single_port_ram11_data_out_net : std_logic_vector( 256-1 downto 0 );
  signal single_port_ram10_data_out_net : std_logic_vector( 256-1 downto 0 );
  signal single_port_ram4_data_out_net : std_logic_vector( 256-1 downto 0 );
  signal single_port_ram13_data_out_net : std_logic_vector( 256-1 downto 0 );
  signal single_port_ram5_data_out_net : std_logic_vector( 256-1 downto 0 );
  signal mux3_y_net : std_logic_vector( 17-1 downto 0 );
  signal single_port_ram6_data_out_net : std_logic_vector( 256-1 downto 0 );
  signal single_port_ram3_data_out_net : std_logic_vector( 256-1 downto 0 );
  signal mux19_y_net : std_logic_vector( 8-1 downto 0 );
  signal single_port_ram8_data_out_net : std_logic_vector( 256-1 downto 0 );
  signal mux28_y_net : std_logic_vector( 17-1 downto 0 );
  signal single_port_ram15_data_out_net : std_logic_vector( 256-1 downto 0 );
  signal mux31_y_net : std_logic_vector( 17-1 downto 0 );
  signal single_port_ram16_data_out_net : std_logic_vector( 256-1 downto 0 );
  signal single_port_ram7_data_out_net : std_logic_vector( 256-1 downto 0 );
  signal mux32_y_net : std_logic_vector( 17-1 downto 0 );
  signal mux35_y_net : std_logic_vector( 17-1 downto 0 );
  signal mux36_y_net : std_logic_vector( 17-1 downto 0 );
  signal mux40_y_net : std_logic_vector( 17-1 downto 0 );
  signal mux39_y_net : std_logic_vector( 17-1 downto 0 );
  signal mux4_y_net : std_logic_vector( 8-1 downto 0 );
  signal mux47_y_net : std_logic_vector( 17-1 downto 0 );
  signal mux48_y_net : std_logic_vector( 17-1 downto 0 );
  signal mux43_y_net : std_logic_vector( 17-1 downto 0 );
  signal mux44_y_net : std_logic_vector( 17-1 downto 0 );
  signal mux56_y_net : std_logic_vector( 17-1 downto 0 );
  signal mux52_y_net : std_logic_vector( 17-1 downto 0 );
  signal mux55_y_net : std_logic_vector( 17-1 downto 0 );
  signal mux5_y_net : std_logic_vector( 8-1 downto 0 );
  signal mux51_y_net : std_logic_vector( 17-1 downto 0 );
  signal mux57_y_net : std_logic_vector( 8-1 downto 0 );
  signal mux8_y_net : std_logic_vector( 8-1 downto 0 );
  signal mux7_y_net : std_logic_vector( 8-1 downto 0 );
  signal mux6_y_net : std_logic_vector( 8-1 downto 0 );
  signal mux9_y_net : std_logic_vector( 8-1 downto 0 );
begin
  out_even1_re <= mux2_y_net;
  out_odd1_re <= mux29_y_net;
  out_even2_re <= mux33_y_net;
  out_odd2_re <= mux37_y_net;
  out_even3_re <= mux41_y_net;
  out_odd3_re <= mux45_y_net;
  out_even4_re <= mux49_y_net;
  out_odd4_re <= mux53_y_net;
  out_even1_im <= mux27_y_net;
  out_odd1_im <= mux30_y_net;
  out_even2_im <= mux34_y_net;
  out_odd2_im <= mux38_y_net;
  out_even3_im <= mux42_y_net;
  out_odd3_im <= mux46_y_net;
  out_even4_im <= mux50_y_net;
  out_odd4_im <= mux54_y_net;
  out_tvalid <= delay11_q_net_x0;
  cordic_6_0_even_1_m_axis_dout_tdata_imag_net_x0 <= in_even1_im;
  cordic_6_0_even_1_m_axis_dout_tdata_real_net_x0 <= in_even1_re;
  cordic_6_0_odd_1_m_axis_dout_tdata_imag_net_x0 <= in_odd1_im;
  cordic_6_0_odd_1_m_axis_dout_tdata_real_net_x0 <= in_odd1_re;
  cordic_6_0_even_2_m_axis_dout_tdata_imag_net_x0 <= in_even2_im;
  cordic_6_0_even_2_m_axis_dout_tdata_real_net_x0 <= in_even2_re;
  cordic_6_0_odd_2_m_axis_dout_tdata_imag_net_x0 <= in_odd2_im;
  cordic_6_0_odd_2_m_axis_dout_tdata_real_net_x0 <= in_odd2_re;
  cordic_6_0_even_1_m_axis_dout_tdata_imag_net <= in_even3_im;
  cordic_6_0_even_1_m_axis_dout_tdata_real_net <= in_even3_re;
  cordic_6_0_odd_1_m_axis_dout_tdata_imag_net <= in_odd3_im;
  cordic_6_0_odd_1_m_axis_dout_tdata_real_net <= in_odd3_re;
  cordic_6_0_even_2_m_axis_dout_tdata_imag_net <= in_even4_im;
  cordic_6_0_even_2_m_axis_dout_tdata_real_net <= in_even4_re;
  cordic_6_0_odd_2_m_axis_dout_tdata_imag_net <= in_odd4_im;
  cordic_6_0_odd_2_m_axis_dout_tdata_real_net <= in_odd4_re;
  cordic_6_0_even_1_m_axis_dout_tvalid_net <= in_tvalid;
  gin_tl_reset_net <= rst;
  delay2_q_net <= data_0;
  delay3_q_net <= data_1;
  delay4_q_net <= data_2;
  delay5_q_net <= data_3;
  delay7_q_net <= data_4;
  delay9_q_net <= data_5;
  delay10_q_net <= data_6;
  delay11_q_net <= data_7;
  delay12_q_net <= w_addr_x0;
  delay16_q_net <= we;
  clk_net <= clk_1;
  ce_net <= ce_1;
  fifo_delay : entity xil_defaultlib.psb3_0_fifo_delay 
  port map (
    in1 => reinterpret32_output_port_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    out1 => fifo3_dout_net_x13
  );
  fifo_delay1 : entity xil_defaultlib.psb3_0_fifo_delay1 
  port map (
    in1 => reinterpret33_output_port_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    out1 => fifo3_dout_net_x12
  );
  fifo_delay10 : entity xil_defaultlib.psb3_0_fifo_delay10 
  port map (
    in1 => reinterpret42_output_port_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    out1 => fifo3_dout_net_x11
  );
  fifo_delay11 : entity xil_defaultlib.psb3_0_fifo_delay11 
  port map (
    in1 => reinterpret43_output_port_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    out1 => fifo3_dout_net_x14
  );
  fifo_delay12 : entity xil_defaultlib.psb3_0_fifo_delay12 
  port map (
    in1 => reinterpret44_output_port_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    out1 => fifo3_dout_net_x10
  );
  fifo_delay13 : entity xil_defaultlib.psb3_0_fifo_delay13 
  port map (
    in1 => reinterpret45_output_port_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    out1 => fifo3_dout_net_x9
  );
  fifo_delay14 : entity xil_defaultlib.psb3_0_fifo_delay14 
  port map (
    in1 => reinterpret46_output_port_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    out1 => fifo3_dout_net_x8
  );
  fifo_delay15 : entity xil_defaultlib.psb3_0_fifo_delay15 
  port map (
    in1 => reinterpret47_output_port_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    out1 => fifo3_dout_net_x7
  );
  fifo_delay2 : entity xil_defaultlib.psb3_0_fifo_delay2 
  port map (
    in1 => reinterpret34_output_port_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    out1 => fifo3_dout_net_x6
  );
  fifo_delay3 : entity xil_defaultlib.psb3_0_fifo_delay3 
  port map (
    in1 => reinterpret35_output_port_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    out1 => fifo3_dout_net_x5
  );
  fifo_delay4 : entity xil_defaultlib.psb3_0_fifo_delay4 
  port map (
    in1 => reinterpret36_output_port_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    out1 => fifo3_dout_net_x4
  );
  fifo_delay5 : entity xil_defaultlib.psb3_0_fifo_delay5 
  port map (
    in1 => reinterpret37_output_port_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    out1 => fifo3_dout_net_x3
  );
  fifo_delay6 : entity xil_defaultlib.psb3_0_fifo_delay6 
  port map (
    in1 => reinterpret38_output_port_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    out1 => fifo3_dout_net_x2
  );
  fifo_delay7 : entity xil_defaultlib.psb3_0_fifo_delay7 
  port map (
    in1 => reinterpret39_output_port_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    out1 => fifo3_dout_net_x1
  );
  fifo_delay8 : entity xil_defaultlib.psb3_0_fifo_delay8 
  port map (
    in1 => reinterpret40_output_port_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    out1 => fifo3_dout_net_x0
  );
  fifo_delay9 : entity xil_defaultlib.psb3_0_fifo_delay9 
  port map (
    in1 => reinterpret41_output_port_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    out1 => fifo3_dout_net
  );
  imag_slice_0 : entity xil_defaultlib.psb3_0_imag_slice_0 
  port map (
    sel => parallel_sel_0_y_net,
    input => mux1_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    output => mux20_y_net_x14
  );
  imag_slice_1 : entity xil_defaultlib.psb3_0_imag_slice_1 
  port map (
    sel => parallel_sel_1_y_net,
    input => mux20_y_net_x15,
    clk_1 => clk_net,
    ce_1 => ce_net,
    output => mux20_y_net_x13
  );
  imag_slice_2 : entity xil_defaultlib.psb3_0_imag_slice_2 
  port map (
    sel => parallel_sel_2_y_net,
    input => mux21_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    output => mux20_y_net_x12
  );
  imag_slice_3 : entity xil_defaultlib.psb3_0_imag_slice_3 
  port map (
    sel => parallel_sel_3_y_net,
    input => mux22_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    output => mux20_y_net_x11
  );
  imag_slice_4 : entity xil_defaultlib.psb3_0_imag_slice_4 
  port map (
    sel => parallel_sel_4_y_net,
    input => mux23_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    output => mux20_y_net_x10
  );
  imag_slice_5 : entity xil_defaultlib.psb3_0_imag_slice_5 
  port map (
    sel => parallel_sel_5_y_net,
    input => mux24_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    output => mux20_y_net_x9
  );
  imag_slice_6 : entity xil_defaultlib.psb3_0_imag_slice_6 
  port map (
    sel => parallel_sel_6_y_net,
    input => mux25_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    output => mux20_y_net_x8
  );
  imag_slice_7 : entity xil_defaultlib.psb3_0_imag_slice_7 
  port map (
    sel => parallel_sel_7_y_net,
    input => mux26_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    output => mux20_y_net_x7
  );
  real_slice_0 : entity xil_defaultlib.psb3_0_real_slice_0 
  port map (
    sel => parallel_sel_0_y_net,
    input => mux1_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    output => mux20_y_net_x6
  );
  real_slice_1 : entity xil_defaultlib.psb3_0_real_slice_1 
  port map (
    sel => parallel_sel_1_y_net,
    input => mux20_y_net_x15,
    clk_1 => clk_net,
    ce_1 => ce_net,
    output => mux20_y_net_x5
  );
  real_slice_2 : entity xil_defaultlib.psb3_0_real_slice_2 
  port map (
    sel => parallel_sel_2_y_net,
    input => mux21_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    output => mux20_y_net_x4
  );
  real_slice_3 : entity xil_defaultlib.psb3_0_real_slice_3 
  port map (
    sel => parallel_sel_3_y_net,
    input => mux22_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    output => mux20_y_net_x3
  );
  real_slice_4 : entity xil_defaultlib.psb3_0_real_slice_4 
  port map (
    sel => parallel_sel_4_y_net,
    input => mux23_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    output => mux20_y_net_x2
  );
  real_slice_5 : entity xil_defaultlib.psb3_0_real_slice_5 
  port map (
    sel => parallel_sel_5_y_net,
    input => mux24_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    output => mux20_y_net_x1
  );
  real_slice_6 : entity xil_defaultlib.psb3_0_real_slice_6 
  port map (
    sel => parallel_sel_6_y_net,
    input => mux25_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    output => mux20_y_net_x0
  );
  real_slice_7 : entity xil_defaultlib.psb3_0_real_slice_7 
  port map (
    sel => parallel_sel_7_y_net,
    input => mux26_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    output => mux20_y_net
  );
  accumulator : entity xil_defaultlib.sysgen_accum_89af09f600 
  port map (
    clr => '0',
    b => relational1_op_net,
    rst => gin_tl_reset_net,
    en => delay13_q_net,
    clk => clk_net,
    ce => ce_net,
    q => accumulator_q_net
  );
  addsub : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 14,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 17,
    core_name0 => "psb3_0_c_addsub_v12_0_i1",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 17,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 17
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret_output_port_net,
    b => reinterpret1_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  addsub1 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 14,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 17,
    core_name0 => "psb3_0_c_addsub_v12_0_i1",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 17,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 17
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret2_output_port_net,
    b => reinterpret3_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  addsub10 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 14,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 17,
    core_name0 => "psb3_0_c_addsub_v12_0_i1",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 17,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 17
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret20_output_port_net,
    b => reinterpret21_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub10_s_net
  );
  addsub11 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 14,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 17,
    core_name0 => "psb3_0_c_addsub_v12_0_i1",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 17,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 17
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret22_output_port_net,
    b => reinterpret23_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub11_s_net
  );
  addsub12 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 14,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 17,
    core_name0 => "psb3_0_c_addsub_v12_0_i1",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 17,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 17
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret24_output_port_net,
    b => reinterpret25_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub12_s_net
  );
  addsub13 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 14,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 17,
    core_name0 => "psb3_0_c_addsub_v12_0_i1",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 17,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 17
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret26_output_port_net,
    b => reinterpret27_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub13_s_net
  );
  addsub14 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 14,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 17,
    core_name0 => "psb3_0_c_addsub_v12_0_i1",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 17,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 17
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret28_output_port_net,
    b => reinterpret29_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub14_s_net
  );
  addsub15 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 14,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 17,
    core_name0 => "psb3_0_c_addsub_v12_0_i1",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 17,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 17
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret30_output_port_net,
    b => reinterpret31_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub15_s_net
  );
  addsub2 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 14,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 17,
    core_name0 => "psb3_0_c_addsub_v12_0_i1",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 17,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 17
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret4_output_port_net,
    b => reinterpret5_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub2_s_net
  );
  addsub3 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 14,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 17,
    core_name0 => "psb3_0_c_addsub_v12_0_i1",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 17,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 17
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret6_output_port_net,
    b => reinterpret7_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub3_s_net
  );
  addsub4 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 14,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 17,
    core_name0 => "psb3_0_c_addsub_v12_0_i1",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 17,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 17
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret8_output_port_net,
    b => reinterpret9_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub4_s_net
  );
  addsub5 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 14,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 17,
    core_name0 => "psb3_0_c_addsub_v12_0_i1",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 17,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 17
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret10_output_port_net,
    b => reinterpret11_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub5_s_net
  );
  addsub6 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 14,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 17,
    core_name0 => "psb3_0_c_addsub_v12_0_i1",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 17,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 17
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret12_output_port_net,
    b => reinterpret13_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub6_s_net
  );
  addsub7 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 14,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 17,
    core_name0 => "psb3_0_c_addsub_v12_0_i1",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 17,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 17
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret14_output_port_net,
    b => reinterpret15_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub7_s_net
  );
  addsub8 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 14,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 17,
    core_name0 => "psb3_0_c_addsub_v12_0_i1",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 17,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 17
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret16_output_port_net,
    b => reinterpret17_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub8_s_net
  );
  addsub9 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 14,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 17,
    core_name0 => "psb3_0_c_addsub_v12_0_i1",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 17,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 17
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret18_output_port_net,
    b => reinterpret19_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub9_s_net
  );
  bitbasher : entity xil_defaultlib.sysgen_bitbasher_8492d24e1e 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    i => addsub_s_net,
    o => bitbasher_o_net
  );
  bitbasher1 : entity xil_defaultlib.sysgen_bitbasher_8492d24e1e 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    i => addsub1_s_net,
    o => bitbasher1_o_net
  );
  bitbasher10 : entity xil_defaultlib.sysgen_bitbasher_8492d24e1e 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    i => addsub10_s_net,
    o => bitbasher10_o_net
  );
  bitbasher11 : entity xil_defaultlib.sysgen_bitbasher_8492d24e1e 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    i => addsub11_s_net,
    o => bitbasher11_o_net
  );
  bitbasher12 : entity xil_defaultlib.sysgen_bitbasher_8492d24e1e 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    i => addsub12_s_net,
    o => bitbasher12_o_net
  );
  bitbasher13 : entity xil_defaultlib.sysgen_bitbasher_8492d24e1e 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    i => addsub13_s_net,
    o => bitbasher13_o_net
  );
  bitbasher14 : entity xil_defaultlib.sysgen_bitbasher_8492d24e1e 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    i => addsub14_s_net,
    o => bitbasher14_o_net
  );
  bitbasher15 : entity xil_defaultlib.sysgen_bitbasher_8492d24e1e 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    i => addsub15_s_net,
    o => bitbasher15_o_net
  );
  bitbasher2 : entity xil_defaultlib.sysgen_bitbasher_8492d24e1e 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    i => addsub2_s_net,
    o => bitbasher2_o_net
  );
  bitbasher3 : entity xil_defaultlib.sysgen_bitbasher_8492d24e1e 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    i => addsub3_s_net,
    o => bitbasher3_o_net
  );
  bitbasher4 : entity xil_defaultlib.sysgen_bitbasher_8492d24e1e 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    i => addsub4_s_net,
    o => bitbasher4_o_net
  );
  bitbasher5 : entity xil_defaultlib.sysgen_bitbasher_8492d24e1e 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    i => addsub5_s_net,
    o => bitbasher5_o_net
  );
  bitbasher6 : entity xil_defaultlib.sysgen_bitbasher_8492d24e1e 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    i => addsub6_s_net,
    o => bitbasher6_o_net
  );
  bitbasher7 : entity xil_defaultlib.sysgen_bitbasher_8492d24e1e 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    i => addsub7_s_net,
    o => bitbasher7_o_net
  );
  bitbasher8 : entity xil_defaultlib.sysgen_bitbasher_8492d24e1e 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    i => addsub8_s_net,
    o => bitbasher8_o_net
  );
  bitbasher9 : entity xil_defaultlib.sysgen_bitbasher_8492d24e1e 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    i => addsub9_s_net,
    o => bitbasher9_o_net
  );
  concat : entity xil_defaultlib.sysgen_concat_6c8db818fa 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => reinterpret32_output_port_net,
    in1 => reinterpret33_output_port_net,
    in2 => reinterpret34_output_port_net,
    in3 => reinterpret35_output_port_net,
    in4 => reinterpret36_output_port_net,
    in5 => reinterpret37_output_port_net,
    in6 => reinterpret38_output_port_net,
    in7 => reinterpret39_output_port_net,
    in8 => reinterpret40_output_port_net,
    in9 => reinterpret41_output_port_net,
    in10 => reinterpret42_output_port_net,
    in11 => reinterpret43_output_port_net,
    in12 => reinterpret44_output_port_net,
    in13 => reinterpret45_output_port_net,
    in14 => reinterpret46_output_port_net,
    in15 => reinterpret47_output_port_net,
    y => concat_y_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_1f1817b2fc 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_f35e175189 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  constant10 : entity xil_defaultlib.sysgen_constant_120ea26d4d 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant10_op_net
  );
  constant11 : entity xil_defaultlib.sysgen_constant_1f1817b2fc 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant11_op_net
  );
  constant12 : entity xil_defaultlib.sysgen_constant_80295d4fb4 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant12_op_net
  );
  constant13 : entity xil_defaultlib.sysgen_constant_1f1817b2fc 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant13_op_net
  );
  constant14 : entity xil_defaultlib.sysgen_constant_e8768a3813 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant14_op_net
  );
  constant15 : entity xil_defaultlib.sysgen_constant_1f1817b2fc 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant15_op_net
  );
  constant16 : entity xil_defaultlib.sysgen_constant_563cb584b0 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant16_op_net
  );
  constant2 : entity xil_defaultlib.sysgen_constant_0714509e7f 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant2_op_net
  );
  constant3 : entity xil_defaultlib.sysgen_constant_1f1817b2fc 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant3_op_net
  );
  constant4 : entity xil_defaultlib.sysgen_constant_754a175f5f 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant4_op_net
  );
  constant5 : entity xil_defaultlib.sysgen_constant_1f1817b2fc 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant5_op_net
  );
  constant6 : entity xil_defaultlib.sysgen_constant_7b0eee2833 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant6_op_net
  );
  constant7 : entity xil_defaultlib.sysgen_constant_1f1817b2fc 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant7_op_net
  );
  constant8 : entity xil_defaultlib.sysgen_constant_d46f498b3d 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant8_op_net
  );
  constant9 : entity xil_defaultlib.sysgen_constant_1f1817b2fc 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant9_op_net
  );
  convert : entity xil_defaultlib.psb3_0_xlconvert 
  generic map (
    bool_conversion => 1,
    din_arith => 1,
    din_bin_pt => 0,
    din_width => 1,
    dout_arith => 1,
    dout_bin_pt => 0,
    dout_width => 1,
    latency => 0,
    overflow => xlWrap,
    quantization => xlTruncate
  )
  port map (
    clr => '0',
    en => "1",
    din => accumulator_q_net,
    clk => clk_net,
    ce => ce_net,
    dout => convert_dout_net
  );
  counter1 : entity xil_defaultlib.psb3_0_xlcounter_free 
  generic map (
    core_name0 => "psb3_0_c_counter_binary_v12_0_i3",
    op_arith => xlUnsigned,
    op_width => 8
  )
  port map (
    clr => '0',
    rst => gin_tl_reset_net,
    en(0) => cordic_6_0_even_1_m_axis_dout_tvalid_net,
    clk => clk_net,
    ce => ce_net,
    op => counter1_op_net
  );
  delay1 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => single_port_ram17_data_out_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay10 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay14_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay10_q_net_x0
  );
  delay11 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 266,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d(0) => cordic_6_0_even_1_m_axis_dout_tvalid_net,
    clk => clk_net,
    ce => ce_net,
    q => delay11_q_net_x0
  );
  delay12 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 4,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => bypass_bool_0_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay12_q_net_x0
  );
  delay13 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 5,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d(0) => cordic_6_0_even_1_m_axis_dout_tvalid_net,
    clk => clk_net,
    ce => ce_net,
    q => delay13_q_net
  );
  delay14 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => convert_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => delay14_q_net
  );
  delay15 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 8
  )
  port map (
    en => '1',
    rst => '0',
    d => counter1_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay15_q_net
  );
  delay16 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 5,
    reg_retiming => 0,
    reset => 0,
    width => 8
  )
  port map (
    en => '1',
    rst => '0',
    d => counter1_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay16_q_net_x0
  );
  delay17 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 8
  )
  port map (
    en => '1',
    rst => '0',
    d => addr_0_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay17_q_net
  );
  delay18 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 4,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => bypass_bool_1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay18_q_net
  );
  delay19 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 5,
    reg_retiming => 0,
    reset => 0,
    width => 8
  )
  port map (
    en => '1',
    rst => '0',
    d => counter1_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay19_q_net
  );
  delay2 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 256
  )
  port map (
    en => '1',
    rst => '0',
    d => concat_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net_x0
  );
  delay20 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 8
  )
  port map (
    en => '1',
    rst => '0',
    d => addr_1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay20_q_net
  );
  delay21 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 4,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => bypass_bool_2_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay21_q_net
  );
  delay22 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 5,
    reg_retiming => 0,
    reset => 0,
    width => 8
  )
  port map (
    en => '1',
    rst => '0',
    d => counter1_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay22_q_net
  );
  delay23 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 8
  )
  port map (
    en => '1',
    rst => '0',
    d => addr_2_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay23_q_net
  );
  delay24 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 4,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => bypass_bool_3_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay24_q_net
  );
  delay25 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 5,
    reg_retiming => 0,
    reset => 0,
    width => 8
  )
  port map (
    en => '1',
    rst => '0',
    d => counter1_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay25_q_net
  );
  delay26 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 8
  )
  port map (
    en => '1',
    rst => '0',
    d => addr_3_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay26_q_net
  );
  delay27 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 4,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => bypass_bool_4_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay27_q_net
  );
  delay28 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 5,
    reg_retiming => 0,
    reset => 0,
    width => 8
  )
  port map (
    en => '1',
    rst => '0',
    d => counter1_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay28_q_net
  );
  delay29 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 8
  )
  port map (
    en => '1',
    rst => '0',
    d => addr_4_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay29_q_net
  );
  delay3 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => single_port_ram18_data_out_net,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net_x0
  );
  delay30 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 4,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => bypass_bool_5_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay30_q_net
  );
  delay31 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 5,
    reg_retiming => 0,
    reset => 0,
    width => 8
  )
  port map (
    en => '1',
    rst => '0',
    d => counter1_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay31_q_net
  );
  delay32 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 8
  )
  port map (
    en => '1',
    rst => '0',
    d => addr_5_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay32_q_net
  );
  delay33 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 4,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => bypass_bool_6_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay33_q_net
  );
  delay34 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 5,
    reg_retiming => 0,
    reset => 0,
    width => 8
  )
  port map (
    en => '1',
    rst => '0',
    d => counter1_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay34_q_net
  );
  delay35 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 8
  )
  port map (
    en => '1',
    rst => '0',
    d => addr_6_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay35_q_net
  );
  delay36 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 4,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => bypass_bool_7_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay36_q_net
  );
  delay37 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 5,
    reg_retiming => 0,
    reset => 0,
    width => 8
  )
  port map (
    en => '1',
    rst => '0',
    d => counter1_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay37_q_net
  );
  delay38 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 8
  )
  port map (
    en => '1',
    rst => '0',
    d => addr_7_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay38_q_net
  );
  delay39 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay16_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay39_q_net
  );
  delay4 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => single_port_ram19_data_out_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net_x0
  );
  delay5 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => single_port_ram20_data_out_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net_x0
  );
  delay6 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => single_port_ram21_data_out_net,
    clk => clk_net,
    ce => ce_net,
    q => delay6_q_net
  );
  delay7 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => single_port_ram22_data_out_net,
    clk => clk_net,
    ce => ce_net,
    q => delay7_q_net_x0
  );
  delay8 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => single_port_ram23_data_out_net,
    clk => clk_net,
    ce => ce_net,
    q => delay8_q_net
  );
  delay9 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => single_port_ram24_data_out_net,
    clk => clk_net,
    ce => ce_net,
    q => delay9_q_net_x0
  );
  inverter : entity xil_defaultlib.sysgen_inverter_ac5174c184 
  port map (
    clr => '0',
    ip => convert_dout_net,
    clk => clk_net,
    ce => ce_net,
    op => inverter_op_net
  );
  logical : entity xil_defaultlib.sysgen_logical_d81059826d 
  port map (
    clr => '0',
    d0 => relational2_op_net,
    d1 => relational_op_net,
    clk => clk_net,
    ce => ce_net,
    y => logical_y_net
  );
  logical1 : entity xil_defaultlib.sysgen_logical_d81059826d 
  port map (
    clr => '0',
    d0 => relational4_op_net,
    d1 => relational3_op_net,
    clk => clk_net,
    ce => ce_net,
    y => logical1_y_net
  );
  logical2 : entity xil_defaultlib.sysgen_logical_d81059826d 
  port map (
    clr => '0',
    d0 => relational6_op_net,
    d1 => relational5_op_net,
    clk => clk_net,
    ce => ce_net,
    y => logical2_y_net
  );
  logical3 : entity xil_defaultlib.sysgen_logical_d81059826d 
  port map (
    clr => '0',
    d0 => relational8_op_net,
    d1 => relational7_op_net,
    clk => clk_net,
    ce => ce_net,
    y => logical3_y_net
  );
  logical4 : entity xil_defaultlib.sysgen_logical_d81059826d 
  port map (
    clr => '0',
    d0 => relational10_op_net,
    d1 => relational9_op_net,
    clk => clk_net,
    ce => ce_net,
    y => logical4_y_net
  );
  logical5 : entity xil_defaultlib.sysgen_logical_d81059826d 
  port map (
    clr => '0',
    d0 => relational12_op_net,
    d1 => relational11_op_net,
    clk => clk_net,
    ce => ce_net,
    y => logical5_y_net
  );
  logical6 : entity xil_defaultlib.sysgen_logical_d81059826d 
  port map (
    clr => '0',
    d0 => relational14_op_net,
    d1 => relational13_op_net,
    clk => clk_net,
    ce => ce_net,
    y => logical6_y_net
  );
  logical7 : entity xil_defaultlib.sysgen_logical_d81059826d 
  port map (
    clr => '0',
    d0 => relational16_op_net,
    d1 => relational15_op_net,
    clk => clk_net,
    ce => ce_net,
    y => logical7_y_net
  );
  mux1 : entity xil_defaultlib.sysgen_mux_1f606cf16b 
  port map (
    clr => '0',
    sel => delay10_q_net_x0,
    d0 => single_port_ram1_data_out_net,
    d1 => single_port_ram9_data_out_net,
    clk => clk_net,
    ce => ce_net,
    y => mux1_y_net
  );
  mux10 : entity xil_defaultlib.sysgen_mux_525d88d897 
  port map (
    clr => '0',
    sel => convert_dout_net,
    d0 => addr_6_y_net,
    d1 => delay15_q_net,
    clk => clk_net,
    ce => ce_net,
    y => mux10_y_net
  );
  mux11 : entity xil_defaultlib.sysgen_mux_525d88d897 
  port map (
    clr => '0',
    sel => convert_dout_net,
    d0 => addr_7_y_net,
    d1 => delay15_q_net,
    clk => clk_net,
    ce => ce_net,
    y => mux11_y_net
  );
  mux12 : entity xil_defaultlib.sysgen_mux_525d88d897 
  port map (
    clr => '0',
    sel => convert_dout_net,
    d0 => delay15_q_net,
    d1 => addr_0_y_net,
    clk => clk_net,
    ce => ce_net,
    y => mux12_y_net
  );
  mux13 : entity xil_defaultlib.sysgen_mux_525d88d897 
  port map (
    clr => '0',
    sel => convert_dout_net,
    d0 => delay15_q_net,
    d1 => addr_1_y_net,
    clk => clk_net,
    ce => ce_net,
    y => mux13_y_net
  );
  mux14 : entity xil_defaultlib.sysgen_mux_525d88d897 
  port map (
    clr => '0',
    sel => convert_dout_net,
    d0 => delay15_q_net,
    d1 => addr_2_y_net,
    clk => clk_net,
    ce => ce_net,
    y => mux14_y_net
  );
  mux15 : entity xil_defaultlib.sysgen_mux_525d88d897 
  port map (
    clr => '0',
    sel => convert_dout_net,
    d0 => delay15_q_net,
    d1 => addr_3_y_net,
    clk => clk_net,
    ce => ce_net,
    y => mux15_y_net
  );
  mux16 : entity xil_defaultlib.sysgen_mux_525d88d897 
  port map (
    clr => '0',
    sel => convert_dout_net,
    d0 => delay15_q_net,
    d1 => addr_4_y_net,
    clk => clk_net,
    ce => ce_net,
    y => mux16_y_net
  );
  mux17 : entity xil_defaultlib.sysgen_mux_525d88d897 
  port map (
    clr => '0',
    sel => convert_dout_net,
    d0 => delay15_q_net,
    d1 => addr_5_y_net,
    clk => clk_net,
    ce => ce_net,
    y => mux17_y_net
  );
  mux18 : entity xil_defaultlib.sysgen_mux_525d88d897 
  port map (
    clr => '0',
    sel => convert_dout_net,
    d0 => delay15_q_net,
    d1 => addr_6_y_net,
    clk => clk_net,
    ce => ce_net,
    y => mux18_y_net
  );
  mux19 : entity xil_defaultlib.sysgen_mux_525d88d897 
  port map (
    clr => '0',
    sel => convert_dout_net,
    d0 => delay15_q_net,
    d1 => addr_7_y_net,
    clk => clk_net,
    ce => ce_net,
    y => mux19_y_net
  );
  mux2 : entity xil_defaultlib.sysgen_mux_32147df3f9 
  port map (
    clr => '0',
    sel => delay12_q_net_x0,
    d0 => constant_op_net,
    d1 => mux3_y_net,
    clk => clk_net,
    ce => ce_net,
    y => mux2_y_net
  );
  mux20 : entity xil_defaultlib.sysgen_mux_1f606cf16b 
  port map (
    clr => '0',
    sel => delay10_q_net_x0,
    d0 => single_port_ram2_data_out_net,
    d1 => single_port_ram10_data_out_net,
    clk => clk_net,
    ce => ce_net,
    y => mux20_y_net_x15
  );
  mux21 : entity xil_defaultlib.sysgen_mux_1f606cf16b 
  port map (
    clr => '0',
    sel => delay10_q_net_x0,
    d0 => single_port_ram3_data_out_net,
    d1 => single_port_ram11_data_out_net,
    clk => clk_net,
    ce => ce_net,
    y => mux21_y_net
  );
  mux22 : entity xil_defaultlib.sysgen_mux_1f606cf16b 
  port map (
    clr => '0',
    sel => delay10_q_net_x0,
    d0 => single_port_ram4_data_out_net,
    d1 => single_port_ram12_data_out_net,
    clk => clk_net,
    ce => ce_net,
    y => mux22_y_net
  );
  mux23 : entity xil_defaultlib.sysgen_mux_1f606cf16b 
  port map (
    clr => '0',
    sel => delay10_q_net_x0,
    d0 => single_port_ram5_data_out_net,
    d1 => single_port_ram13_data_out_net,
    clk => clk_net,
    ce => ce_net,
    y => mux23_y_net
  );
  mux24 : entity xil_defaultlib.sysgen_mux_1f606cf16b 
  port map (
    clr => '0',
    sel => delay10_q_net_x0,
    d0 => single_port_ram6_data_out_net,
    d1 => single_port_ram14_data_out_net,
    clk => clk_net,
    ce => ce_net,
    y => mux24_y_net
  );
  mux25 : entity xil_defaultlib.sysgen_mux_1f606cf16b 
  port map (
    clr => '0',
    sel => delay10_q_net_x0,
    d0 => single_port_ram7_data_out_net,
    d1 => single_port_ram15_data_out_net,
    clk => clk_net,
    ce => ce_net,
    y => mux25_y_net
  );
  mux26 : entity xil_defaultlib.sysgen_mux_1f606cf16b 
  port map (
    clr => '0',
    sel => delay10_q_net_x0,
    d0 => single_port_ram8_data_out_net,
    d1 => single_port_ram16_data_out_net,
    clk => clk_net,
    ce => ce_net,
    y => mux26_y_net
  );
  mux27 : entity xil_defaultlib.sysgen_mux_32147df3f9 
  port map (
    clr => '0',
    sel => delay12_q_net_x0,
    d0 => constant_op_net,
    d1 => mux28_y_net,
    clk => clk_net,
    ce => ce_net,
    y => mux27_y_net
  );
  mux28 : entity xil_defaultlib.sysgen_mux_32147df3f9 
  port map (
    clr => '0',
    sel => logical_y_net,
    d0 => addsub1_s_net,
    d1 => bitbasher1_o_net,
    clk => clk_net,
    ce => ce_net,
    y => mux28_y_net
  );
  mux29 : entity xil_defaultlib.sysgen_mux_32147df3f9 
  port map (
    clr => '0',
    sel => delay18_q_net,
    d0 => constant3_op_net,
    d1 => mux32_y_net,
    clk => clk_net,
    ce => ce_net,
    y => mux29_y_net
  );
  mux3 : entity xil_defaultlib.sysgen_mux_32147df3f9 
  port map (
    clr => '0',
    sel => logical_y_net,
    d0 => addsub_s_net,
    d1 => bitbasher_o_net,
    clk => clk_net,
    ce => ce_net,
    y => mux3_y_net
  );
  mux30 : entity xil_defaultlib.sysgen_mux_32147df3f9 
  port map (
    clr => '0',
    sel => delay18_q_net,
    d0 => constant3_op_net,
    d1 => mux31_y_net,
    clk => clk_net,
    ce => ce_net,
    y => mux30_y_net
  );
  mux31 : entity xil_defaultlib.sysgen_mux_32147df3f9 
  port map (
    clr => '0',
    sel => logical1_y_net,
    d0 => addsub3_s_net,
    d1 => bitbasher3_o_net,
    clk => clk_net,
    ce => ce_net,
    y => mux31_y_net
  );
  mux32 : entity xil_defaultlib.sysgen_mux_32147df3f9 
  port map (
    clr => '0',
    sel => logical1_y_net,
    d0 => addsub2_s_net,
    d1 => bitbasher2_o_net,
    clk => clk_net,
    ce => ce_net,
    y => mux32_y_net
  );
  mux33 : entity xil_defaultlib.sysgen_mux_32147df3f9 
  port map (
    clr => '0',
    sel => delay21_q_net,
    d0 => constant5_op_net,
    d1 => mux36_y_net,
    clk => clk_net,
    ce => ce_net,
    y => mux33_y_net
  );
  mux34 : entity xil_defaultlib.sysgen_mux_32147df3f9 
  port map (
    clr => '0',
    sel => delay21_q_net,
    d0 => constant5_op_net,
    d1 => mux35_y_net,
    clk => clk_net,
    ce => ce_net,
    y => mux34_y_net
  );
  mux35 : entity xil_defaultlib.sysgen_mux_32147df3f9 
  port map (
    clr => '0',
    sel => logical2_y_net,
    d0 => addsub5_s_net,
    d1 => bitbasher5_o_net,
    clk => clk_net,
    ce => ce_net,
    y => mux35_y_net
  );
  mux36 : entity xil_defaultlib.sysgen_mux_32147df3f9 
  port map (
    clr => '0',
    sel => logical2_y_net,
    d0 => addsub4_s_net,
    d1 => bitbasher4_o_net,
    clk => clk_net,
    ce => ce_net,
    y => mux36_y_net
  );
  mux37 : entity xil_defaultlib.sysgen_mux_32147df3f9 
  port map (
    clr => '0',
    sel => delay24_q_net,
    d0 => constant7_op_net,
    d1 => mux40_y_net,
    clk => clk_net,
    ce => ce_net,
    y => mux37_y_net
  );
  mux38 : entity xil_defaultlib.sysgen_mux_32147df3f9 
  port map (
    clr => '0',
    sel => delay24_q_net,
    d0 => constant7_op_net,
    d1 => mux39_y_net,
    clk => clk_net,
    ce => ce_net,
    y => mux38_y_net
  );
  mux39 : entity xil_defaultlib.sysgen_mux_32147df3f9 
  port map (
    clr => '0',
    sel => logical3_y_net,
    d0 => addsub7_s_net,
    d1 => bitbasher7_o_net,
    clk => clk_net,
    ce => ce_net,
    y => mux39_y_net
  );
  mux4 : entity xil_defaultlib.sysgen_mux_525d88d897 
  port map (
    clr => '0',
    sel => convert_dout_net,
    d0 => addr_0_y_net,
    d1 => delay15_q_net,
    clk => clk_net,
    ce => ce_net,
    y => mux4_y_net
  );
  mux40 : entity xil_defaultlib.sysgen_mux_32147df3f9 
  port map (
    clr => '0',
    sel => logical3_y_net,
    d0 => addsub6_s_net,
    d1 => bitbasher6_o_net,
    clk => clk_net,
    ce => ce_net,
    y => mux40_y_net
  );
  mux41 : entity xil_defaultlib.sysgen_mux_32147df3f9 
  port map (
    clr => '0',
    sel => delay27_q_net,
    d0 => constant9_op_net,
    d1 => mux44_y_net,
    clk => clk_net,
    ce => ce_net,
    y => mux41_y_net
  );
  mux42 : entity xil_defaultlib.sysgen_mux_32147df3f9 
  port map (
    clr => '0',
    sel => delay27_q_net,
    d0 => constant9_op_net,
    d1 => mux43_y_net,
    clk => clk_net,
    ce => ce_net,
    y => mux42_y_net
  );
  mux43 : entity xil_defaultlib.sysgen_mux_32147df3f9 
  port map (
    clr => '0',
    sel => logical4_y_net,
    d0 => addsub9_s_net,
    d1 => bitbasher9_o_net,
    clk => clk_net,
    ce => ce_net,
    y => mux43_y_net
  );
  mux44 : entity xil_defaultlib.sysgen_mux_32147df3f9 
  port map (
    clr => '0',
    sel => logical4_y_net,
    d0 => addsub8_s_net,
    d1 => bitbasher8_o_net,
    clk => clk_net,
    ce => ce_net,
    y => mux44_y_net
  );
  mux45 : entity xil_defaultlib.sysgen_mux_32147df3f9 
  port map (
    clr => '0',
    sel => delay30_q_net,
    d0 => constant11_op_net,
    d1 => mux48_y_net,
    clk => clk_net,
    ce => ce_net,
    y => mux45_y_net
  );
  mux46 : entity xil_defaultlib.sysgen_mux_32147df3f9 
  port map (
    clr => '0',
    sel => delay30_q_net,
    d0 => constant11_op_net,
    d1 => mux47_y_net,
    clk => clk_net,
    ce => ce_net,
    y => mux46_y_net
  );
  mux47 : entity xil_defaultlib.sysgen_mux_32147df3f9 
  port map (
    clr => '0',
    sel => logical5_y_net,
    d0 => addsub11_s_net,
    d1 => bitbasher11_o_net,
    clk => clk_net,
    ce => ce_net,
    y => mux47_y_net
  );
  mux48 : entity xil_defaultlib.sysgen_mux_32147df3f9 
  port map (
    clr => '0',
    sel => logical5_y_net,
    d0 => addsub10_s_net,
    d1 => bitbasher10_o_net,
    clk => clk_net,
    ce => ce_net,
    y => mux48_y_net
  );
  mux49 : entity xil_defaultlib.sysgen_mux_32147df3f9 
  port map (
    clr => '0',
    sel => delay33_q_net,
    d0 => constant13_op_net,
    d1 => mux52_y_net,
    clk => clk_net,
    ce => ce_net,
    y => mux49_y_net
  );
  mux5 : entity xil_defaultlib.sysgen_mux_525d88d897 
  port map (
    clr => '0',
    sel => convert_dout_net,
    d0 => addr_1_y_net,
    d1 => delay15_q_net,
    clk => clk_net,
    ce => ce_net,
    y => mux5_y_net
  );
  mux50 : entity xil_defaultlib.sysgen_mux_32147df3f9 
  port map (
    clr => '0',
    sel => delay33_q_net,
    d0 => constant13_op_net,
    d1 => mux51_y_net,
    clk => clk_net,
    ce => ce_net,
    y => mux50_y_net
  );
  mux51 : entity xil_defaultlib.sysgen_mux_32147df3f9 
  port map (
    clr => '0',
    sel => logical6_y_net,
    d0 => addsub13_s_net,
    d1 => bitbasher13_o_net,
    clk => clk_net,
    ce => ce_net,
    y => mux51_y_net
  );
  mux52 : entity xil_defaultlib.sysgen_mux_32147df3f9 
  port map (
    clr => '0',
    sel => logical6_y_net,
    d0 => addsub12_s_net,
    d1 => bitbasher12_o_net,
    clk => clk_net,
    ce => ce_net,
    y => mux52_y_net
  );
  mux53 : entity xil_defaultlib.sysgen_mux_32147df3f9 
  port map (
    clr => '0',
    sel => delay36_q_net,
    d0 => constant15_op_net,
    d1 => mux56_y_net,
    clk => clk_net,
    ce => ce_net,
    y => mux53_y_net
  );
  mux54 : entity xil_defaultlib.sysgen_mux_32147df3f9 
  port map (
    clr => '0',
    sel => delay36_q_net,
    d0 => constant15_op_net,
    d1 => mux55_y_net,
    clk => clk_net,
    ce => ce_net,
    y => mux54_y_net
  );
  mux55 : entity xil_defaultlib.sysgen_mux_32147df3f9 
  port map (
    clr => '0',
    sel => logical7_y_net,
    d0 => addsub15_s_net,
    d1 => bitbasher15_o_net,
    clk => clk_net,
    ce => ce_net,
    y => mux55_y_net
  );
  mux56 : entity xil_defaultlib.sysgen_mux_32147df3f9 
  port map (
    clr => '0',
    sel => logical7_y_net,
    d0 => addsub14_s_net,
    d1 => bitbasher14_o_net,
    clk => clk_net,
    ce => ce_net,
    y => mux56_y_net
  );
  mux57 : entity xil_defaultlib.sysgen_mux_525d88d897 
  port map (
    clr => '0',
    sel => delay16_q_net,
    d0 => counter1_op_net,
    d1 => delay12_q_net,
    clk => clk_net,
    ce => ce_net,
    y => mux57_y_net
  );
  mux6 : entity xil_defaultlib.sysgen_mux_525d88d897 
  port map (
    clr => '0',
    sel => convert_dout_net,
    d0 => addr_2_y_net,
    d1 => delay15_q_net,
    clk => clk_net,
    ce => ce_net,
    y => mux6_y_net
  );
  mux7 : entity xil_defaultlib.sysgen_mux_525d88d897 
  port map (
    clr => '0',
    sel => convert_dout_net,
    d0 => addr_3_y_net,
    d1 => delay15_q_net,
    clk => clk_net,
    ce => ce_net,
    y => mux7_y_net
  );
  mux8 : entity xil_defaultlib.sysgen_mux_525d88d897 
  port map (
    clr => '0',
    sel => convert_dout_net,
    d0 => addr_4_y_net,
    d1 => delay15_q_net,
    clk => clk_net,
    ce => ce_net,
    y => mux8_y_net
  );
  mux9 : entity xil_defaultlib.sysgen_mux_525d88d897 
  port map (
    clr => '0',
    sel => convert_dout_net,
    d0 => addr_5_y_net,
    d1 => delay15_q_net,
    clk => clk_net,
    ce => ce_net,
    y => mux9_y_net
  );
  reinterpret : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => fifo3_dout_net_x7,
    output_port => reinterpret_output_port_net
  );
  reinterpret1 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => mux20_y_net_x6,
    output_port => reinterpret1_output_port_net
  );
  reinterpret10 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => fifo3_dout_net_x11,
    output_port => reinterpret10_output_port_net
  );
  reinterpret11 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => mux20_y_net_x12,
    output_port => reinterpret11_output_port_net
  );
  reinterpret12 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => fifo3_dout_net,
    output_port => reinterpret12_output_port_net
  );
  reinterpret13 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => mux20_y_net_x3,
    output_port => reinterpret13_output_port_net
  );
  reinterpret14 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => fifo3_dout_net_x0,
    output_port => reinterpret14_output_port_net
  );
  reinterpret15 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => mux20_y_net_x11,
    output_port => reinterpret15_output_port_net
  );
  reinterpret16 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => fifo3_dout_net_x1,
    output_port => reinterpret16_output_port_net
  );
  reinterpret17 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => mux20_y_net_x2,
    output_port => reinterpret17_output_port_net
  );
  reinterpret18 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => fifo3_dout_net_x2,
    output_port => reinterpret18_output_port_net
  );
  reinterpret19 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => mux20_y_net_x10,
    output_port => reinterpret19_output_port_net
  );
  reinterpret2 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => fifo3_dout_net_x8,
    output_port => reinterpret2_output_port_net
  );
  reinterpret20 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => fifo3_dout_net_x3,
    output_port => reinterpret20_output_port_net
  );
  reinterpret21 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => mux20_y_net_x1,
    output_port => reinterpret21_output_port_net
  );
  reinterpret22 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => fifo3_dout_net_x4,
    output_port => reinterpret22_output_port_net
  );
  reinterpret23 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => mux20_y_net_x9,
    output_port => reinterpret23_output_port_net
  );
  reinterpret24 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => fifo3_dout_net_x5,
    output_port => reinterpret24_output_port_net
  );
  reinterpret25 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => mux20_y_net_x0,
    output_port => reinterpret25_output_port_net
  );
  reinterpret26 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => fifo3_dout_net_x6,
    output_port => reinterpret26_output_port_net
  );
  reinterpret27 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => mux20_y_net_x8,
    output_port => reinterpret27_output_port_net
  );
  reinterpret28 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => fifo3_dout_net_x12,
    output_port => reinterpret28_output_port_net
  );
  reinterpret29 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => mux20_y_net,
    output_port => reinterpret29_output_port_net
  );
  reinterpret3 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => mux20_y_net_x14,
    output_port => reinterpret3_output_port_net
  );
  reinterpret30 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => fifo3_dout_net_x13,
    output_port => reinterpret30_output_port_net
  );
  reinterpret31 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => mux20_y_net_x7,
    output_port => reinterpret31_output_port_net
  );
  reinterpret32 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => cordic_6_0_odd_2_m_axis_dout_tdata_imag_net,
    output_port => reinterpret32_output_port_net
  );
  reinterpret33 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => cordic_6_0_odd_2_m_axis_dout_tdata_real_net,
    output_port => reinterpret33_output_port_net
  );
  reinterpret34 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => cordic_6_0_even_2_m_axis_dout_tdata_imag_net,
    output_port => reinterpret34_output_port_net
  );
  reinterpret35 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => cordic_6_0_even_2_m_axis_dout_tdata_real_net,
    output_port => reinterpret35_output_port_net
  );
  reinterpret36 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => cordic_6_0_odd_1_m_axis_dout_tdata_imag_net,
    output_port => reinterpret36_output_port_net
  );
  reinterpret37 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => cordic_6_0_odd_1_m_axis_dout_tdata_real_net,
    output_port => reinterpret37_output_port_net
  );
  reinterpret38 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => cordic_6_0_even_1_m_axis_dout_tdata_imag_net,
    output_port => reinterpret38_output_port_net
  );
  reinterpret39 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => cordic_6_0_even_1_m_axis_dout_tdata_real_net,
    output_port => reinterpret39_output_port_net
  );
  reinterpret4 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => fifo3_dout_net_x9,
    output_port => reinterpret4_output_port_net
  );
  reinterpret40 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => cordic_6_0_odd_2_m_axis_dout_tdata_imag_net_x0,
    output_port => reinterpret40_output_port_net
  );
  reinterpret41 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => cordic_6_0_odd_2_m_axis_dout_tdata_real_net_x0,
    output_port => reinterpret41_output_port_net
  );
  reinterpret42 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => cordic_6_0_even_2_m_axis_dout_tdata_imag_net_x0,
    output_port => reinterpret42_output_port_net
  );
  reinterpret43 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => cordic_6_0_even_2_m_axis_dout_tdata_real_net_x0,
    output_port => reinterpret43_output_port_net
  );
  reinterpret44 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => cordic_6_0_odd_1_m_axis_dout_tdata_imag_net_x0,
    output_port => reinterpret44_output_port_net
  );
  reinterpret45 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => cordic_6_0_odd_1_m_axis_dout_tdata_real_net_x0,
    output_port => reinterpret45_output_port_net
  );
  reinterpret46 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => cordic_6_0_even_1_m_axis_dout_tdata_imag_net_x0,
    output_port => reinterpret46_output_port_net
  );
  reinterpret47 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => cordic_6_0_even_1_m_axis_dout_tdata_real_net_x0,
    output_port => reinterpret47_output_port_net
  );
  reinterpret5 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => mux20_y_net_x5,
    output_port => reinterpret5_output_port_net
  );
  reinterpret6 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => fifo3_dout_net_x10,
    output_port => reinterpret6_output_port_net
  );
  reinterpret7 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => mux20_y_net_x13,
    output_port => reinterpret7_output_port_net
  );
  reinterpret8 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => fifo3_dout_net_x14,
    output_port => reinterpret8_output_port_net
  );
  reinterpret9 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => mux20_y_net_x4,
    output_port => reinterpret9_output_port_net
  );
  relational : entity xil_defaultlib.sysgen_relational_5aa8d67ef0 
  port map (
    clr => '0',
    a => constant1_op_net,
    b => parallel_sel_0_y_net,
    clk => clk_net,
    ce => ce_net,
    op => relational_op_net
  );
  relational1 : entity xil_defaultlib.sysgen_relational_226ad2322f 
  port map (
    clr => '0',
    a => counter1_op_net,
    b => constant2_op_net,
    clk => clk_net,
    ce => ce_net,
    op => relational1_op_net
  );
  relational10 : entity xil_defaultlib.sysgen_relational_d1682fb355 
  port map (
    clr => '0',
    a => delay28_q_net,
    b => delay29_q_net,
    clk => clk_net,
    ce => ce_net,
    op => relational10_op_net
  );
  relational11 : entity xil_defaultlib.sysgen_relational_5aa8d67ef0 
  port map (
    clr => '0',
    a => constant12_op_net,
    b => parallel_sel_5_y_net,
    clk => clk_net,
    ce => ce_net,
    op => relational11_op_net
  );
  relational12 : entity xil_defaultlib.sysgen_relational_d1682fb355 
  port map (
    clr => '0',
    a => delay31_q_net,
    b => delay32_q_net,
    clk => clk_net,
    ce => ce_net,
    op => relational12_op_net
  );
  relational13 : entity xil_defaultlib.sysgen_relational_5aa8d67ef0 
  port map (
    clr => '0',
    a => constant14_op_net,
    b => parallel_sel_6_y_net,
    clk => clk_net,
    ce => ce_net,
    op => relational13_op_net
  );
  relational14 : entity xil_defaultlib.sysgen_relational_d1682fb355 
  port map (
    clr => '0',
    a => delay34_q_net,
    b => delay35_q_net,
    clk => clk_net,
    ce => ce_net,
    op => relational14_op_net
  );
  relational15 : entity xil_defaultlib.sysgen_relational_5aa8d67ef0 
  port map (
    clr => '0',
    a => constant16_op_net,
    b => parallel_sel_7_y_net,
    clk => clk_net,
    ce => ce_net,
    op => relational15_op_net
  );
  relational16 : entity xil_defaultlib.sysgen_relational_d1682fb355 
  port map (
    clr => '0',
    a => delay37_q_net,
    b => delay38_q_net,
    clk => clk_net,
    ce => ce_net,
    op => relational16_op_net
  );
  relational2 : entity xil_defaultlib.sysgen_relational_d1682fb355 
  port map (
    clr => '0',
    a => delay16_q_net_x0,
    b => delay17_q_net,
    clk => clk_net,
    ce => ce_net,
    op => relational2_op_net
  );
  relational3 : entity xil_defaultlib.sysgen_relational_5aa8d67ef0 
  port map (
    clr => '0',
    a => constant4_op_net,
    b => parallel_sel_1_y_net,
    clk => clk_net,
    ce => ce_net,
    op => relational3_op_net
  );
  relational4 : entity xil_defaultlib.sysgen_relational_d1682fb355 
  port map (
    clr => '0',
    a => delay19_q_net,
    b => delay20_q_net,
    clk => clk_net,
    ce => ce_net,
    op => relational4_op_net
  );
  relational5 : entity xil_defaultlib.sysgen_relational_5aa8d67ef0 
  port map (
    clr => '0',
    a => constant6_op_net,
    b => parallel_sel_2_y_net,
    clk => clk_net,
    ce => ce_net,
    op => relational5_op_net
  );
  relational6 : entity xil_defaultlib.sysgen_relational_d1682fb355 
  port map (
    clr => '0',
    a => delay22_q_net,
    b => delay23_q_net,
    clk => clk_net,
    ce => ce_net,
    op => relational6_op_net
  );
  relational7 : entity xil_defaultlib.sysgen_relational_5aa8d67ef0 
  port map (
    clr => '0',
    a => constant8_op_net,
    b => parallel_sel_3_y_net,
    clk => clk_net,
    ce => ce_net,
    op => relational7_op_net
  );
  relational8 : entity xil_defaultlib.sysgen_relational_d1682fb355 
  port map (
    clr => '0',
    a => delay25_q_net,
    b => delay26_q_net,
    clk => clk_net,
    ce => ce_net,
    op => relational8_op_net
  );
  relational9 : entity xil_defaultlib.sysgen_relational_5aa8d67ef0 
  port map (
    clr => '0',
    a => constant10_op_net,
    b => parallel_sel_4_y_net,
    clk => clk_net,
    ce => ce_net,
    op => relational9_op_net
  );
  single_port_ram1 : entity xil_defaultlib.psb3_0_xlspram 
  generic map (
    init_value => b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
    latency => 1,
    mem_init_file => "xpm_4dd9cf_vivado.mem",
    mem_size => 65536,
    mem_type => "block",
    read_reset_val => "0",
    width => 256,
    width_addr => 8,
    write_mode_a => "write_first",
    xpm_lat => 1
  )
  port map (
    en => "1",
    rst => "0",
    addr => mux4_y_net,
    data_in => delay2_q_net_x0,
    we => delay14_q_net,
    clk => clk_net,
    ce => ce_net,
    data_out => single_port_ram1_data_out_net
  );
  single_port_ram10 : entity xil_defaultlib.psb3_0_xlspram 
  generic map (
    init_value => b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
    latency => 1,
    mem_init_file => "xpm_4dd9cf_vivado.mem",
    mem_size => 65536,
    mem_type => "block",
    read_reset_val => "0",
    width => 256,
    width_addr => 8,
    write_mode_a => "write_first",
    xpm_lat => 1
  )
  port map (
    en => "1",
    rst => "0",
    addr => mux13_y_net,
    data_in => delay2_q_net_x0,
    we => inverter_op_net,
    clk => clk_net,
    ce => ce_net,
    data_out => single_port_ram10_data_out_net
  );
  single_port_ram11 : entity xil_defaultlib.psb3_0_xlspram 
  generic map (
    init_value => b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
    latency => 1,
    mem_init_file => "xpm_4dd9cf_vivado.mem",
    mem_size => 65536,
    mem_type => "block",
    read_reset_val => "0",
    width => 256,
    width_addr => 8,
    write_mode_a => "write_first",
    xpm_lat => 1
  )
  port map (
    en => "1",
    rst => "0",
    addr => mux14_y_net,
    data_in => delay2_q_net_x0,
    we => inverter_op_net,
    clk => clk_net,
    ce => ce_net,
    data_out => single_port_ram11_data_out_net
  );
  single_port_ram12 : entity xil_defaultlib.psb3_0_xlspram 
  generic map (
    init_value => b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
    latency => 1,
    mem_init_file => "xpm_4dd9cf_vivado.mem",
    mem_size => 65536,
    mem_type => "block",
    read_reset_val => "0",
    width => 256,
    width_addr => 8,
    write_mode_a => "write_first",
    xpm_lat => 1
  )
  port map (
    en => "1",
    rst => "0",
    addr => mux15_y_net,
    data_in => delay2_q_net_x0,
    we => inverter_op_net,
    clk => clk_net,
    ce => ce_net,
    data_out => single_port_ram12_data_out_net
  );
  single_port_ram13 : entity xil_defaultlib.psb3_0_xlspram 
  generic map (
    init_value => b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
    latency => 1,
    mem_init_file => "xpm_4dd9cf_vivado.mem",
    mem_size => 65536,
    mem_type => "block",
    read_reset_val => "0",
    width => 256,
    width_addr => 8,
    write_mode_a => "write_first",
    xpm_lat => 1
  )
  port map (
    en => "1",
    rst => "0",
    addr => mux16_y_net,
    data_in => delay2_q_net_x0,
    we => inverter_op_net,
    clk => clk_net,
    ce => ce_net,
    data_out => single_port_ram13_data_out_net
  );
  single_port_ram14 : entity xil_defaultlib.psb3_0_xlspram 
  generic map (
    init_value => b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
    latency => 1,
    mem_init_file => "xpm_4dd9cf_vivado.mem",
    mem_size => 65536,
    mem_type => "block",
    read_reset_val => "0",
    width => 256,
    width_addr => 8,
    write_mode_a => "write_first",
    xpm_lat => 1
  )
  port map (
    en => "1",
    rst => "0",
    addr => mux17_y_net,
    data_in => delay2_q_net_x0,
    we => inverter_op_net,
    clk => clk_net,
    ce => ce_net,
    data_out => single_port_ram14_data_out_net
  );
  single_port_ram15 : entity xil_defaultlib.psb3_0_xlspram 
  generic map (
    init_value => b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
    latency => 1,
    mem_init_file => "xpm_4dd9cf_vivado.mem",
    mem_size => 65536,
    mem_type => "block",
    read_reset_val => "0",
    width => 256,
    width_addr => 8,
    write_mode_a => "write_first",
    xpm_lat => 1
  )
  port map (
    en => "1",
    rst => "0",
    addr => mux18_y_net,
    data_in => delay2_q_net_x0,
    we => inverter_op_net,
    clk => clk_net,
    ce => ce_net,
    data_out => single_port_ram15_data_out_net
  );
  single_port_ram16 : entity xil_defaultlib.psb3_0_xlspram 
  generic map (
    init_value => b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
    latency => 1,
    mem_init_file => "xpm_4dd9cf_vivado.mem",
    mem_size => 65536,
    mem_type => "block",
    read_reset_val => "0",
    width => 256,
    width_addr => 8,
    write_mode_a => "write_first",
    xpm_lat => 1
  )
  port map (
    en => "1",
    rst => "0",
    addr => mux19_y_net,
    data_in => delay2_q_net_x0,
    we => inverter_op_net,
    clk => clk_net,
    ce => ce_net,
    data_out => single_port_ram16_data_out_net
  );
  single_port_ram17 : entity xil_defaultlib.psb3_0_xlspram 
  generic map (
    init_value => b"000000000000",
    latency => 1,
    mem_init_file => "xpm_763daf_vivado.mem",
    mem_size => 3072,
    mem_type => "block",
    read_reset_val => "0",
    width => 12,
    width_addr => 8,
    write_mode_a => "write_first",
    xpm_lat => 1
  )
  port map (
    en => "1",
    rst => "0",
    addr => mux57_y_net,
    data_in => delay2_q_net,
    we => delay39_q_net,
    clk => clk_net,
    ce => ce_net,
    data_out => single_port_ram17_data_out_net
  );
  single_port_ram18 : entity xil_defaultlib.psb3_0_xlspram 
  generic map (
    init_value => b"000000000000",
    latency => 1,
    mem_init_file => "xpm_5ecc77_vivado.mem",
    mem_size => 3072,
    mem_type => "block",
    read_reset_val => "0",
    width => 12,
    width_addr => 8,
    write_mode_a => "write_first",
    xpm_lat => 1
  )
  port map (
    en => "1",
    rst => "0",
    addr => mux57_y_net,
    data_in => delay3_q_net,
    we => delay39_q_net,
    clk => clk_net,
    ce => ce_net,
    data_out => single_port_ram18_data_out_net
  );
  single_port_ram19 : entity xil_defaultlib.psb3_0_xlspram 
  generic map (
    init_value => b"000000000000",
    latency => 1,
    mem_init_file => "xpm_5c779c_vivado.mem",
    mem_size => 3072,
    mem_type => "block",
    read_reset_val => "0",
    width => 12,
    width_addr => 8,
    write_mode_a => "write_first",
    xpm_lat => 1
  )
  port map (
    en => "1",
    rst => "0",
    addr => mux57_y_net,
    data_in => delay4_q_net,
    we => delay39_q_net,
    clk => clk_net,
    ce => ce_net,
    data_out => single_port_ram19_data_out_net
  );
  single_port_ram2 : entity xil_defaultlib.psb3_0_xlspram 
  generic map (
    init_value => b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
    latency => 1,
    mem_init_file => "xpm_4dd9cf_vivado.mem",
    mem_size => 65536,
    mem_type => "block",
    read_reset_val => "0",
    width => 256,
    width_addr => 8,
    write_mode_a => "write_first",
    xpm_lat => 1
  )
  port map (
    en => "1",
    rst => "0",
    addr => mux5_y_net,
    data_in => delay2_q_net_x0,
    we => delay14_q_net,
    clk => clk_net,
    ce => ce_net,
    data_out => single_port_ram2_data_out_net
  );
  single_port_ram20 : entity xil_defaultlib.psb3_0_xlspram 
  generic map (
    init_value => b"000000000000",
    latency => 1,
    mem_init_file => "xpm_1937ca_vivado.mem",
    mem_size => 3072,
    mem_type => "block",
    read_reset_val => "0",
    width => 12,
    width_addr => 8,
    write_mode_a => "write_first",
    xpm_lat => 1
  )
  port map (
    en => "1",
    rst => "0",
    addr => mux57_y_net,
    data_in => delay5_q_net,
    we => delay39_q_net,
    clk => clk_net,
    ce => ce_net,
    data_out => single_port_ram20_data_out_net
  );
  single_port_ram21 : entity xil_defaultlib.psb3_0_xlspram 
  generic map (
    init_value => b"000000000000",
    latency => 1,
    mem_init_file => "xpm_af1f98_vivado.mem",
    mem_size => 3072,
    mem_type => "block",
    read_reset_val => "0",
    width => 12,
    width_addr => 8,
    write_mode_a => "write_first",
    xpm_lat => 1
  )
  port map (
    en => "1",
    rst => "0",
    addr => mux57_y_net,
    data_in => delay7_q_net,
    we => delay39_q_net,
    clk => clk_net,
    ce => ce_net,
    data_out => single_port_ram21_data_out_net
  );
  single_port_ram22 : entity xil_defaultlib.psb3_0_xlspram 
  generic map (
    init_value => b"000000000000",
    latency => 1,
    mem_init_file => "xpm_4b85a4_vivado.mem",
    mem_size => 3072,
    mem_type => "block",
    read_reset_val => "0",
    width => 12,
    width_addr => 8,
    write_mode_a => "write_first",
    xpm_lat => 1
  )
  port map (
    en => "1",
    rst => "0",
    addr => mux57_y_net,
    data_in => delay9_q_net,
    we => delay39_q_net,
    clk => clk_net,
    ce => ce_net,
    data_out => single_port_ram22_data_out_net
  );
  single_port_ram23 : entity xil_defaultlib.psb3_0_xlspram 
  generic map (
    init_value => b"000000000000",
    latency => 1,
    mem_init_file => "xpm_ff0e07_vivado.mem",
    mem_size => 3072,
    mem_type => "block",
    read_reset_val => "0",
    width => 12,
    width_addr => 8,
    write_mode_a => "write_first",
    xpm_lat => 1
  )
  port map (
    en => "1",
    rst => "0",
    addr => mux57_y_net,
    data_in => delay10_q_net,
    we => delay39_q_net,
    clk => clk_net,
    ce => ce_net,
    data_out => single_port_ram23_data_out_net
  );
  single_port_ram24 : entity xil_defaultlib.psb3_0_xlspram 
  generic map (
    init_value => b"000000000000",
    latency => 1,
    mem_init_file => "xpm_7bf015_vivado.mem",
    mem_size => 3072,
    mem_type => "block",
    read_reset_val => "0",
    width => 12,
    width_addr => 8,
    write_mode_a => "write_first",
    xpm_lat => 1
  )
  port map (
    en => "1",
    rst => "0",
    addr => mux57_y_net,
    data_in => delay11_q_net,
    we => delay39_q_net,
    clk => clk_net,
    ce => ce_net,
    data_out => single_port_ram24_data_out_net
  );
  single_port_ram3 : entity xil_defaultlib.psb3_0_xlspram 
  generic map (
    init_value => b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
    latency => 1,
    mem_init_file => "xpm_4dd9cf_vivado.mem",
    mem_size => 65536,
    mem_type => "block",
    read_reset_val => "0",
    width => 256,
    width_addr => 8,
    write_mode_a => "write_first",
    xpm_lat => 1
  )
  port map (
    en => "1",
    rst => "0",
    addr => mux6_y_net,
    data_in => delay2_q_net_x0,
    we => delay14_q_net,
    clk => clk_net,
    ce => ce_net,
    data_out => single_port_ram3_data_out_net
  );
  single_port_ram4 : entity xil_defaultlib.psb3_0_xlspram 
  generic map (
    init_value => b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
    latency => 1,
    mem_init_file => "xpm_4dd9cf_vivado.mem",
    mem_size => 65536,
    mem_type => "block",
    read_reset_val => "0",
    width => 256,
    width_addr => 8,
    write_mode_a => "write_first",
    xpm_lat => 1
  )
  port map (
    en => "1",
    rst => "0",
    addr => mux7_y_net,
    data_in => delay2_q_net_x0,
    we => delay14_q_net,
    clk => clk_net,
    ce => ce_net,
    data_out => single_port_ram4_data_out_net
  );
  single_port_ram5 : entity xil_defaultlib.psb3_0_xlspram 
  generic map (
    init_value => b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
    latency => 1,
    mem_init_file => "xpm_4dd9cf_vivado.mem",
    mem_size => 65536,
    mem_type => "block",
    read_reset_val => "0",
    width => 256,
    width_addr => 8,
    write_mode_a => "write_first",
    xpm_lat => 1
  )
  port map (
    en => "1",
    rst => "0",
    addr => mux8_y_net,
    data_in => delay2_q_net_x0,
    we => delay14_q_net,
    clk => clk_net,
    ce => ce_net,
    data_out => single_port_ram5_data_out_net
  );
  single_port_ram6 : entity xil_defaultlib.psb3_0_xlspram 
  generic map (
    init_value => b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
    latency => 1,
    mem_init_file => "xpm_4dd9cf_vivado.mem",
    mem_size => 65536,
    mem_type => "block",
    read_reset_val => "0",
    width => 256,
    width_addr => 8,
    write_mode_a => "write_first",
    xpm_lat => 1
  )
  port map (
    en => "1",
    rst => "0",
    addr => mux9_y_net,
    data_in => delay2_q_net_x0,
    we => delay14_q_net,
    clk => clk_net,
    ce => ce_net,
    data_out => single_port_ram6_data_out_net
  );
  single_port_ram7 : entity xil_defaultlib.psb3_0_xlspram 
  generic map (
    init_value => b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
    latency => 1,
    mem_init_file => "xpm_4dd9cf_vivado.mem",
    mem_size => 65536,
    mem_type => "block",
    read_reset_val => "0",
    width => 256,
    width_addr => 8,
    write_mode_a => "write_first",
    xpm_lat => 1
  )
  port map (
    en => "1",
    rst => "0",
    addr => mux10_y_net,
    data_in => delay2_q_net_x0,
    we => delay14_q_net,
    clk => clk_net,
    ce => ce_net,
    data_out => single_port_ram7_data_out_net
  );
  single_port_ram8 : entity xil_defaultlib.psb3_0_xlspram 
  generic map (
    init_value => b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
    latency => 1,
    mem_init_file => "xpm_4dd9cf_vivado.mem",
    mem_size => 65536,
    mem_type => "block",
    read_reset_val => "0",
    width => 256,
    width_addr => 8,
    write_mode_a => "write_first",
    xpm_lat => 1
  )
  port map (
    en => "1",
    rst => "0",
    addr => mux11_y_net,
    data_in => delay2_q_net_x0,
    we => delay14_q_net,
    clk => clk_net,
    ce => ce_net,
    data_out => single_port_ram8_data_out_net
  );
  single_port_ram9 : entity xil_defaultlib.psb3_0_xlspram 
  generic map (
    init_value => b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
    latency => 1,
    mem_init_file => "xpm_4dd9cf_vivado.mem",
    mem_size => 65536,
    mem_type => "block",
    read_reset_val => "0",
    width => 256,
    width_addr => 8,
    write_mode_a => "write_first",
    xpm_lat => 1
  )
  port map (
    en => "1",
    rst => "0",
    addr => mux12_y_net,
    data_in => delay2_q_net_x0,
    we => inverter_op_net,
    clk => clk_net,
    ce => ce_net,
    data_out => single_port_ram9_data_out_net
  );
  addr_0 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 4,
    new_msb => 11,
    x_width => 12,
    y_width => 8
  )
  port map (
    x => single_port_ram17_data_out_net,
    y => addr_0_y_net
  );
  addr_1 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 4,
    new_msb => 11,
    x_width => 12,
    y_width => 8
  )
  port map (
    x => single_port_ram18_data_out_net,
    y => addr_1_y_net
  );
  addr_2 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 4,
    new_msb => 11,
    x_width => 12,
    y_width => 8
  )
  port map (
    x => single_port_ram19_data_out_net,
    y => addr_2_y_net
  );
  addr_3 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 4,
    new_msb => 11,
    x_width => 12,
    y_width => 8
  )
  port map (
    x => single_port_ram20_data_out_net,
    y => addr_3_y_net
  );
  addr_4 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 4,
    new_msb => 11,
    x_width => 12,
    y_width => 8
  )
  port map (
    x => single_port_ram21_data_out_net,
    y => addr_4_y_net
  );
  addr_5 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 4,
    new_msb => 11,
    x_width => 12,
    y_width => 8
  )
  port map (
    x => single_port_ram22_data_out_net,
    y => addr_5_y_net
  );
  addr_6 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 4,
    new_msb => 11,
    x_width => 12,
    y_width => 8
  )
  port map (
    x => single_port_ram23_data_out_net,
    y => addr_6_y_net
  );
  addr_7 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 4,
    new_msb => 11,
    x_width => 12,
    y_width => 8
  )
  port map (
    x => single_port_ram24_data_out_net,
    y => addr_7_y_net
  );
  bypass_bool_0 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 0,
    x_width => 12,
    y_width => 1
  )
  port map (
    x => delay1_q_net,
    y => bypass_bool_0_y_net
  );
  bypass_bool_1 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 0,
    x_width => 12,
    y_width => 1
  )
  port map (
    x => delay3_q_net_x0,
    y => bypass_bool_1_y_net
  );
  bypass_bool_2 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 0,
    x_width => 12,
    y_width => 1
  )
  port map (
    x => delay4_q_net_x0,
    y => bypass_bool_2_y_net
  );
  bypass_bool_3 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 0,
    x_width => 12,
    y_width => 1
  )
  port map (
    x => delay5_q_net_x0,
    y => bypass_bool_3_y_net
  );
  bypass_bool_4 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 0,
    x_width => 12,
    y_width => 1
  )
  port map (
    x => delay6_q_net,
    y => bypass_bool_4_y_net
  );
  bypass_bool_5 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 0,
    x_width => 12,
    y_width => 1
  )
  port map (
    x => delay7_q_net_x0,
    y => bypass_bool_5_y_net
  );
  bypass_bool_6 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 0,
    x_width => 12,
    y_width => 1
  )
  port map (
    x => delay8_q_net,
    y => bypass_bool_6_y_net
  );
  bypass_bool_7 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 0,
    x_width => 12,
    y_width => 1
  )
  port map (
    x => delay9_q_net_x0,
    y => bypass_bool_7_y_net
  );
  parallel_sel_0 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 1,
    new_msb => 3,
    x_width => 12,
    y_width => 3
  )
  port map (
    x => delay1_q_net,
    y => parallel_sel_0_y_net
  );
  parallel_sel_1 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 1,
    new_msb => 3,
    x_width => 12,
    y_width => 3
  )
  port map (
    x => delay3_q_net_x0,
    y => parallel_sel_1_y_net
  );
  parallel_sel_2 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 1,
    new_msb => 3,
    x_width => 12,
    y_width => 3
  )
  port map (
    x => delay4_q_net_x0,
    y => parallel_sel_2_y_net
  );
  parallel_sel_3 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 1,
    new_msb => 3,
    x_width => 12,
    y_width => 3
  )
  port map (
    x => delay5_q_net_x0,
    y => parallel_sel_3_y_net
  );
  parallel_sel_4 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 1,
    new_msb => 3,
    x_width => 12,
    y_width => 3
  )
  port map (
    x => delay6_q_net,
    y => parallel_sel_4_y_net
  );
  parallel_sel_5 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 1,
    new_msb => 3,
    x_width => 12,
    y_width => 3
  )
  port map (
    x => delay7_q_net_x0,
    y => parallel_sel_5_y_net
  );
  parallel_sel_6 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 1,
    new_msb => 3,
    x_width => 12,
    y_width => 3
  )
  port map (
    x => delay8_q_net,
    y => parallel_sel_6_y_net
  );
  parallel_sel_7 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 1,
    new_msb => 3,
    x_width => 12,
    y_width => 3
  )
  port map (
    x => delay9_q_net_x0,
    y => parallel_sel_7_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Vector AddSub Fabric
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_addsub_fabric is
  port (
    a_1 : in std_logic_vector( 16-1 downto 0 );
    b_1 : in std_logic_vector( 16-1 downto 0 );
    a_2 : in std_logic_vector( 16-1 downto 0 );
    a_3 : in std_logic_vector( 16-1 downto 0 );
    a_4 : in std_logic_vector( 16-1 downto 0 );
    a_5 : in std_logic_vector( 16-1 downto 0 );
    a_6 : in std_logic_vector( 16-1 downto 0 );
    a_7 : in std_logic_vector( 16-1 downto 0 );
    a_8 : in std_logic_vector( 16-1 downto 0 );
    a_9 : in std_logic_vector( 16-1 downto 0 );
    a_10 : in std_logic_vector( 16-1 downto 0 );
    a_11 : in std_logic_vector( 16-1 downto 0 );
    a_12 : in std_logic_vector( 16-1 downto 0 );
    a_13 : in std_logic_vector( 16-1 downto 0 );
    a_14 : in std_logic_vector( 16-1 downto 0 );
    a_15 : in std_logic_vector( 16-1 downto 0 );
    a_16 : in std_logic_vector( 16-1 downto 0 );
    b_2 : in std_logic_vector( 16-1 downto 0 );
    b_3 : in std_logic_vector( 16-1 downto 0 );
    b_4 : in std_logic_vector( 16-1 downto 0 );
    b_5 : in std_logic_vector( 16-1 downto 0 );
    b_6 : in std_logic_vector( 16-1 downto 0 );
    b_7 : in std_logic_vector( 16-1 downto 0 );
    b_8 : in std_logic_vector( 16-1 downto 0 );
    b_9 : in std_logic_vector( 16-1 downto 0 );
    b_10 : in std_logic_vector( 16-1 downto 0 );
    b_11 : in std_logic_vector( 16-1 downto 0 );
    b_12 : in std_logic_vector( 16-1 downto 0 );
    b_13 : in std_logic_vector( 16-1 downto 0 );
    b_14 : in std_logic_vector( 16-1 downto 0 );
    b_15 : in std_logic_vector( 16-1 downto 0 );
    b_16 : in std_logic_vector( 16-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    a_b_1 : out std_logic_vector( 16-1 downto 0 );
    a_b_2 : out std_logic_vector( 16-1 downto 0 );
    a_b_3 : out std_logic_vector( 16-1 downto 0 );
    a_b_4 : out std_logic_vector( 16-1 downto 0 );
    a_b_5 : out std_logic_vector( 16-1 downto 0 );
    a_b_6 : out std_logic_vector( 16-1 downto 0 );
    a_b_7 : out std_logic_vector( 16-1 downto 0 );
    a_b_8 : out std_logic_vector( 16-1 downto 0 );
    a_b_9 : out std_logic_vector( 16-1 downto 0 );
    a_b_10 : out std_logic_vector( 16-1 downto 0 );
    a_b_11 : out std_logic_vector( 16-1 downto 0 );
    a_b_12 : out std_logic_vector( 16-1 downto 0 );
    a_b_13 : out std_logic_vector( 16-1 downto 0 );
    a_b_14 : out std_logic_vector( 16-1 downto 0 );
    a_b_15 : out std_logic_vector( 16-1 downto 0 );
    a_b_16 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_vector_addsub_fabric;
architecture structural of psb3_0_vector_addsub_fabric is 
  signal addsub0_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub5_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub3_s_net : std_logic_vector( 16-1 downto 0 );
  signal mult4_p_net : std_logic_vector( 16-1 downto 0 );
  signal addsub15_s_net : std_logic_vector( 16-1 downto 0 );
  signal mult9_p_net : std_logic_vector( 16-1 downto 0 );
  signal addsub10_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub12_s_net : std_logic_vector( 16-1 downto 0 );
  signal mult2_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult0_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult1_p_net : std_logic_vector( 16-1 downto 0 );
  signal addsub11_s_net : std_logic_vector( 16-1 downto 0 );
  signal mult3_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult8_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult12_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult13_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult5_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult10_p_net : std_logic_vector( 16-1 downto 0 );
  signal addsub7_s_net : std_logic_vector( 16-1 downto 0 );
  signal mult6_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult7_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult14_p_net : std_logic_vector( 16-1 downto 0 );
  signal addsub14_s_net : std_logic_vector( 16-1 downto 0 );
  signal mult15_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub9_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub8_s_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mult11_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub13_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub6_s_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal clk_net : std_logic;
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal ce_net : std_logic;
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
begin
  a_b_1 <= addsub0_s_net;
  a_b_2 <= addsub1_s_net;
  a_b_3 <= addsub2_s_net;
  a_b_4 <= addsub3_s_net;
  a_b_5 <= addsub4_s_net;
  a_b_6 <= addsub5_s_net;
  a_b_7 <= addsub6_s_net;
  a_b_8 <= addsub7_s_net;
  a_b_9 <= addsub8_s_net;
  a_b_10 <= addsub9_s_net;
  a_b_11 <= addsub10_s_net;
  a_b_12 <= addsub11_s_net;
  a_b_13 <= addsub12_s_net;
  a_b_14 <= addsub13_s_net;
  a_b_15 <= addsub14_s_net;
  a_b_16 <= addsub15_s_net;
  mult0_p_net <= a_1;
  reinterpret0_output_port_net <= b_1;
  mult1_p_net <= a_2;
  mult2_p_net <= a_3;
  mult3_p_net <= a_4;
  mult4_p_net <= a_5;
  mult5_p_net <= a_6;
  mult6_p_net <= a_7;
  mult7_p_net <= a_8;
  mult8_p_net <= a_9;
  mult9_p_net <= a_10;
  mult10_p_net <= a_11;
  mult11_p_net <= a_12;
  mult12_p_net <= a_13;
  mult13_p_net <= a_14;
  mult14_p_net <= a_15;
  mult15_p_net <= a_16;
  reinterpret1_output_port_net <= b_2;
  reinterpret2_output_port_net <= b_3;
  reinterpret3_output_port_net <= b_4;
  reinterpret4_output_port_net <= b_5;
  reinterpret5_output_port_net <= b_6;
  reinterpret6_output_port_net <= b_7;
  reinterpret7_output_port_net <= b_8;
  reinterpret8_output_port_net <= b_9;
  reinterpret9_output_port_net <= b_10;
  reinterpret10_output_port_net <= b_11;
  reinterpret11_output_port_net <= b_12;
  reinterpret12_output_port_net <= b_13;
  reinterpret13_output_port_net <= b_14;
  reinterpret14_output_port_net <= b_15;
  reinterpret15_output_port_net <= b_16;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub0 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult0_p_net,
    b => reinterpret0_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub0_s_net
  );
  addsub1 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult1_p_net,
    b => reinterpret1_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  addsub2 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult2_p_net,
    b => reinterpret2_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub2_s_net
  );
  addsub3 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult3_p_net,
    b => reinterpret3_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub3_s_net
  );
  addsub4 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult4_p_net,
    b => reinterpret4_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub4_s_net
  );
  addsub5 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult5_p_net,
    b => reinterpret5_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub5_s_net
  );
  addsub6 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult6_p_net,
    b => reinterpret6_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub6_s_net
  );
  addsub7 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult7_p_net,
    b => reinterpret7_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub7_s_net
  );
  addsub8 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult8_p_net,
    b => reinterpret8_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub8_s_net
  );
  addsub9 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult9_p_net,
    b => reinterpret9_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub9_s_net
  );
  addsub10 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult10_p_net,
    b => reinterpret10_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub10_s_net
  );
  addsub11 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult11_p_net,
    b => reinterpret11_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub11_s_net
  );
  addsub12 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult12_p_net,
    b => reinterpret12_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub12_s_net
  );
  addsub13 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult13_p_net,
    b => reinterpret13_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub13_s_net
  );
  addsub14 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult14_p_net,
    b => reinterpret14_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub14_s_net
  );
  addsub15 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult15_p_net,
    b => reinterpret15_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub15_s_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Vector AddSub Fabric1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_addsub_fabric1 is
  port (
    a_1 : in std_logic_vector( 16-1 downto 0 );
    b_1 : in std_logic_vector( 16-1 downto 0 );
    a_2 : in std_logic_vector( 16-1 downto 0 );
    a_3 : in std_logic_vector( 16-1 downto 0 );
    a_4 : in std_logic_vector( 16-1 downto 0 );
    a_5 : in std_logic_vector( 16-1 downto 0 );
    a_6 : in std_logic_vector( 16-1 downto 0 );
    a_7 : in std_logic_vector( 16-1 downto 0 );
    a_8 : in std_logic_vector( 16-1 downto 0 );
    a_9 : in std_logic_vector( 16-1 downto 0 );
    a_10 : in std_logic_vector( 16-1 downto 0 );
    a_11 : in std_logic_vector( 16-1 downto 0 );
    a_12 : in std_logic_vector( 16-1 downto 0 );
    a_13 : in std_logic_vector( 16-1 downto 0 );
    a_14 : in std_logic_vector( 16-1 downto 0 );
    a_15 : in std_logic_vector( 16-1 downto 0 );
    a_16 : in std_logic_vector( 16-1 downto 0 );
    b_2 : in std_logic_vector( 16-1 downto 0 );
    b_3 : in std_logic_vector( 16-1 downto 0 );
    b_4 : in std_logic_vector( 16-1 downto 0 );
    b_5 : in std_logic_vector( 16-1 downto 0 );
    b_6 : in std_logic_vector( 16-1 downto 0 );
    b_7 : in std_logic_vector( 16-1 downto 0 );
    b_8 : in std_logic_vector( 16-1 downto 0 );
    b_9 : in std_logic_vector( 16-1 downto 0 );
    b_10 : in std_logic_vector( 16-1 downto 0 );
    b_11 : in std_logic_vector( 16-1 downto 0 );
    b_12 : in std_logic_vector( 16-1 downto 0 );
    b_13 : in std_logic_vector( 16-1 downto 0 );
    b_14 : in std_logic_vector( 16-1 downto 0 );
    b_15 : in std_logic_vector( 16-1 downto 0 );
    b_16 : in std_logic_vector( 16-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    a_b_1 : out std_logic_vector( 16-1 downto 0 );
    a_b_2 : out std_logic_vector( 16-1 downto 0 );
    a_b_3 : out std_logic_vector( 16-1 downto 0 );
    a_b_4 : out std_logic_vector( 16-1 downto 0 );
    a_b_5 : out std_logic_vector( 16-1 downto 0 );
    a_b_6 : out std_logic_vector( 16-1 downto 0 );
    a_b_7 : out std_logic_vector( 16-1 downto 0 );
    a_b_8 : out std_logic_vector( 16-1 downto 0 );
    a_b_9 : out std_logic_vector( 16-1 downto 0 );
    a_b_10 : out std_logic_vector( 16-1 downto 0 );
    a_b_11 : out std_logic_vector( 16-1 downto 0 );
    a_b_12 : out std_logic_vector( 16-1 downto 0 );
    a_b_13 : out std_logic_vector( 16-1 downto 0 );
    a_b_14 : out std_logic_vector( 16-1 downto 0 );
    a_b_15 : out std_logic_vector( 16-1 downto 0 );
    a_b_16 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_vector_addsub_fabric1;
architecture structural of psb3_0_vector_addsub_fabric1 is 
  signal mult9_p_net : std_logic_vector( 16-1 downto 0 );
  signal addsub12_s_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mult2_p_net : std_logic_vector( 16-1 downto 0 );
  signal addsub3_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub5_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub10_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 16-1 downto 0 );
  signal mult1_p_net : std_logic_vector( 16-1 downto 0 );
  signal addsub6_s_net : std_logic_vector( 16-1 downto 0 );
  signal mult3_p_net : std_logic_vector( 16-1 downto 0 );
  signal addsub7_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub9_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub11_s_net : std_logic_vector( 16-1 downto 0 );
  signal mult0_p_net : std_logic_vector( 16-1 downto 0 );
  signal addsub14_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub13_s_net : std_logic_vector( 16-1 downto 0 );
  signal mult4_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult5_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult6_p_net : std_logic_vector( 16-1 downto 0 );
  signal addsub15_s_net : std_logic_vector( 16-1 downto 0 );
  signal mult7_p_net : std_logic_vector( 16-1 downto 0 );
  signal addsub0_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub8_s_net : std_logic_vector( 16-1 downto 0 );
  signal mult8_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal clk_net : std_logic;
  signal ce_net : std_logic;
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mult10_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult14_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mult15_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult13_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult11_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult12_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
begin
  a_b_1 <= addsub0_s_net;
  a_b_2 <= addsub1_s_net;
  a_b_3 <= addsub2_s_net;
  a_b_4 <= addsub3_s_net;
  a_b_5 <= addsub4_s_net;
  a_b_6 <= addsub5_s_net;
  a_b_7 <= addsub6_s_net;
  a_b_8 <= addsub7_s_net;
  a_b_9 <= addsub8_s_net;
  a_b_10 <= addsub9_s_net;
  a_b_11 <= addsub10_s_net;
  a_b_12 <= addsub11_s_net;
  a_b_13 <= addsub12_s_net;
  a_b_14 <= addsub13_s_net;
  a_b_15 <= addsub14_s_net;
  a_b_16 <= addsub15_s_net;
  mult0_p_net <= a_1;
  reinterpret0_output_port_net <= b_1;
  mult1_p_net <= a_2;
  mult2_p_net <= a_3;
  mult3_p_net <= a_4;
  mult4_p_net <= a_5;
  mult5_p_net <= a_6;
  mult6_p_net <= a_7;
  mult7_p_net <= a_8;
  mult8_p_net <= a_9;
  mult9_p_net <= a_10;
  mult10_p_net <= a_11;
  mult11_p_net <= a_12;
  mult12_p_net <= a_13;
  mult13_p_net <= a_14;
  mult14_p_net <= a_15;
  mult15_p_net <= a_16;
  reinterpret1_output_port_net <= b_2;
  reinterpret2_output_port_net <= b_3;
  reinterpret3_output_port_net <= b_4;
  reinterpret4_output_port_net <= b_5;
  reinterpret5_output_port_net <= b_6;
  reinterpret6_output_port_net <= b_7;
  reinterpret7_output_port_net <= b_8;
  reinterpret8_output_port_net <= b_9;
  reinterpret9_output_port_net <= b_10;
  reinterpret10_output_port_net <= b_11;
  reinterpret11_output_port_net <= b_12;
  reinterpret12_output_port_net <= b_13;
  reinterpret13_output_port_net <= b_14;
  reinterpret14_output_port_net <= b_15;
  reinterpret15_output_port_net <= b_16;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub0 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult0_p_net,
    b => reinterpret0_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub0_s_net
  );
  addsub1 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult1_p_net,
    b => reinterpret1_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  addsub2 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult2_p_net,
    b => reinterpret2_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub2_s_net
  );
  addsub3 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult3_p_net,
    b => reinterpret3_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub3_s_net
  );
  addsub4 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult4_p_net,
    b => reinterpret4_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub4_s_net
  );
  addsub5 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult5_p_net,
    b => reinterpret5_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub5_s_net
  );
  addsub6 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult6_p_net,
    b => reinterpret6_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub6_s_net
  );
  addsub7 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult7_p_net,
    b => reinterpret7_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub7_s_net
  );
  addsub8 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult8_p_net,
    b => reinterpret8_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub8_s_net
  );
  addsub9 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult9_p_net,
    b => reinterpret9_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub9_s_net
  );
  addsub10 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult10_p_net,
    b => reinterpret10_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub10_s_net
  );
  addsub11 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult11_p_net,
    b => reinterpret11_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub11_s_net
  );
  addsub12 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult12_p_net,
    b => reinterpret12_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub12_s_net
  );
  addsub13 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult13_p_net,
    b => reinterpret13_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub13_s_net
  );
  addsub14 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult14_p_net,
    b => reinterpret14_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub14_s_net
  );
  addsub15 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult15_p_net,
    b => reinterpret15_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub15_s_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Vector AddSub Fabric2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_addsub_fabric2 is
  port (
    a_1 : in std_logic_vector( 16-1 downto 0 );
    b_1 : in std_logic_vector( 16-1 downto 0 );
    a_2 : in std_logic_vector( 16-1 downto 0 );
    a_3 : in std_logic_vector( 16-1 downto 0 );
    a_4 : in std_logic_vector( 16-1 downto 0 );
    a_5 : in std_logic_vector( 16-1 downto 0 );
    a_6 : in std_logic_vector( 16-1 downto 0 );
    a_7 : in std_logic_vector( 16-1 downto 0 );
    a_8 : in std_logic_vector( 16-1 downto 0 );
    a_9 : in std_logic_vector( 16-1 downto 0 );
    a_10 : in std_logic_vector( 16-1 downto 0 );
    a_11 : in std_logic_vector( 16-1 downto 0 );
    a_12 : in std_logic_vector( 16-1 downto 0 );
    a_13 : in std_logic_vector( 16-1 downto 0 );
    a_14 : in std_logic_vector( 16-1 downto 0 );
    a_15 : in std_logic_vector( 16-1 downto 0 );
    a_16 : in std_logic_vector( 16-1 downto 0 );
    b_2 : in std_logic_vector( 16-1 downto 0 );
    b_3 : in std_logic_vector( 16-1 downto 0 );
    b_4 : in std_logic_vector( 16-1 downto 0 );
    b_5 : in std_logic_vector( 16-1 downto 0 );
    b_6 : in std_logic_vector( 16-1 downto 0 );
    b_7 : in std_logic_vector( 16-1 downto 0 );
    b_8 : in std_logic_vector( 16-1 downto 0 );
    b_9 : in std_logic_vector( 16-1 downto 0 );
    b_10 : in std_logic_vector( 16-1 downto 0 );
    b_11 : in std_logic_vector( 16-1 downto 0 );
    b_12 : in std_logic_vector( 16-1 downto 0 );
    b_13 : in std_logic_vector( 16-1 downto 0 );
    b_14 : in std_logic_vector( 16-1 downto 0 );
    b_15 : in std_logic_vector( 16-1 downto 0 );
    b_16 : in std_logic_vector( 16-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    a_b_1 : out std_logic_vector( 16-1 downto 0 );
    a_b_2 : out std_logic_vector( 16-1 downto 0 );
    a_b_3 : out std_logic_vector( 16-1 downto 0 );
    a_b_4 : out std_logic_vector( 16-1 downto 0 );
    a_b_5 : out std_logic_vector( 16-1 downto 0 );
    a_b_6 : out std_logic_vector( 16-1 downto 0 );
    a_b_7 : out std_logic_vector( 16-1 downto 0 );
    a_b_8 : out std_logic_vector( 16-1 downto 0 );
    a_b_9 : out std_logic_vector( 16-1 downto 0 );
    a_b_10 : out std_logic_vector( 16-1 downto 0 );
    a_b_11 : out std_logic_vector( 16-1 downto 0 );
    a_b_12 : out std_logic_vector( 16-1 downto 0 );
    a_b_13 : out std_logic_vector( 16-1 downto 0 );
    a_b_14 : out std_logic_vector( 16-1 downto 0 );
    a_b_15 : out std_logic_vector( 16-1 downto 0 );
    a_b_16 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_vector_addsub_fabric2;
architecture structural of psb3_0_vector_addsub_fabric2 is 
  signal addsub4_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub6_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub8_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub9_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub10_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub5_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub12_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub3_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub13_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub14_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub7_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub11_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub15_s_net : std_logic_vector( 16-1 downto 0 );
  signal mult0_p_net : std_logic_vector( 16-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub0_s_net : std_logic_vector( 16-1 downto 0 );
  signal clk_net : std_logic;
  signal mult14_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mult11_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mult4_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult5_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult9_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mult3_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult2_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult15_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mult8_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mult6_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mult13_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult10_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mult7_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult12_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult1_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal ce_net : std_logic;
begin
  a_b_1 <= addsub0_s_net;
  a_b_2 <= addsub1_s_net;
  a_b_3 <= addsub2_s_net;
  a_b_4 <= addsub3_s_net;
  a_b_5 <= addsub4_s_net;
  a_b_6 <= addsub5_s_net;
  a_b_7 <= addsub6_s_net;
  a_b_8 <= addsub7_s_net;
  a_b_9 <= addsub8_s_net;
  a_b_10 <= addsub9_s_net;
  a_b_11 <= addsub10_s_net;
  a_b_12 <= addsub11_s_net;
  a_b_13 <= addsub12_s_net;
  a_b_14 <= addsub13_s_net;
  a_b_15 <= addsub14_s_net;
  a_b_16 <= addsub15_s_net;
  mult0_p_net <= a_1;
  reinterpret0_output_port_net <= b_1;
  mult1_p_net <= a_2;
  mult2_p_net <= a_3;
  mult3_p_net <= a_4;
  mult4_p_net <= a_5;
  mult5_p_net <= a_6;
  mult6_p_net <= a_7;
  mult7_p_net <= a_8;
  mult8_p_net <= a_9;
  mult9_p_net <= a_10;
  mult10_p_net <= a_11;
  mult11_p_net <= a_12;
  mult12_p_net <= a_13;
  mult13_p_net <= a_14;
  mult14_p_net <= a_15;
  mult15_p_net <= a_16;
  reinterpret1_output_port_net <= b_2;
  reinterpret2_output_port_net <= b_3;
  reinterpret3_output_port_net <= b_4;
  reinterpret4_output_port_net <= b_5;
  reinterpret5_output_port_net <= b_6;
  reinterpret6_output_port_net <= b_7;
  reinterpret7_output_port_net <= b_8;
  reinterpret8_output_port_net <= b_9;
  reinterpret9_output_port_net <= b_10;
  reinterpret10_output_port_net <= b_11;
  reinterpret11_output_port_net <= b_12;
  reinterpret12_output_port_net <= b_13;
  reinterpret13_output_port_net <= b_14;
  reinterpret14_output_port_net <= b_15;
  reinterpret15_output_port_net <= b_16;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub0 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult0_p_net,
    b => reinterpret0_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub0_s_net
  );
  addsub1 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult1_p_net,
    b => reinterpret1_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  addsub2 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult2_p_net,
    b => reinterpret2_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub2_s_net
  );
  addsub3 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult3_p_net,
    b => reinterpret3_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub3_s_net
  );
  addsub4 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult4_p_net,
    b => reinterpret4_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub4_s_net
  );
  addsub5 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult5_p_net,
    b => reinterpret5_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub5_s_net
  );
  addsub6 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult6_p_net,
    b => reinterpret6_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub6_s_net
  );
  addsub7 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult7_p_net,
    b => reinterpret7_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub7_s_net
  );
  addsub8 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult8_p_net,
    b => reinterpret8_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub8_s_net
  );
  addsub9 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult9_p_net,
    b => reinterpret9_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub9_s_net
  );
  addsub10 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult10_p_net,
    b => reinterpret10_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub10_s_net
  );
  addsub11 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult11_p_net,
    b => reinterpret11_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub11_s_net
  );
  addsub12 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult12_p_net,
    b => reinterpret12_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub12_s_net
  );
  addsub13 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult13_p_net,
    b => reinterpret13_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub13_s_net
  );
  addsub14 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult14_p_net,
    b => reinterpret14_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub14_s_net
  );
  addsub15 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult15_p_net,
    b => reinterpret15_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub15_s_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Vector AddSub Fabric3
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_addsub_fabric3 is
  port (
    a_1 : in std_logic_vector( 16-1 downto 0 );
    b_1 : in std_logic_vector( 16-1 downto 0 );
    a_2 : in std_logic_vector( 16-1 downto 0 );
    a_3 : in std_logic_vector( 16-1 downto 0 );
    a_4 : in std_logic_vector( 16-1 downto 0 );
    a_5 : in std_logic_vector( 16-1 downto 0 );
    a_6 : in std_logic_vector( 16-1 downto 0 );
    a_7 : in std_logic_vector( 16-1 downto 0 );
    a_8 : in std_logic_vector( 16-1 downto 0 );
    a_9 : in std_logic_vector( 16-1 downto 0 );
    a_10 : in std_logic_vector( 16-1 downto 0 );
    a_11 : in std_logic_vector( 16-1 downto 0 );
    a_12 : in std_logic_vector( 16-1 downto 0 );
    a_13 : in std_logic_vector( 16-1 downto 0 );
    a_14 : in std_logic_vector( 16-1 downto 0 );
    a_15 : in std_logic_vector( 16-1 downto 0 );
    a_16 : in std_logic_vector( 16-1 downto 0 );
    b_2 : in std_logic_vector( 16-1 downto 0 );
    b_3 : in std_logic_vector( 16-1 downto 0 );
    b_4 : in std_logic_vector( 16-1 downto 0 );
    b_5 : in std_logic_vector( 16-1 downto 0 );
    b_6 : in std_logic_vector( 16-1 downto 0 );
    b_7 : in std_logic_vector( 16-1 downto 0 );
    b_8 : in std_logic_vector( 16-1 downto 0 );
    b_9 : in std_logic_vector( 16-1 downto 0 );
    b_10 : in std_logic_vector( 16-1 downto 0 );
    b_11 : in std_logic_vector( 16-1 downto 0 );
    b_12 : in std_logic_vector( 16-1 downto 0 );
    b_13 : in std_logic_vector( 16-1 downto 0 );
    b_14 : in std_logic_vector( 16-1 downto 0 );
    b_15 : in std_logic_vector( 16-1 downto 0 );
    b_16 : in std_logic_vector( 16-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    a_b_1 : out std_logic_vector( 16-1 downto 0 );
    a_b_2 : out std_logic_vector( 16-1 downto 0 );
    a_b_3 : out std_logic_vector( 16-1 downto 0 );
    a_b_4 : out std_logic_vector( 16-1 downto 0 );
    a_b_5 : out std_logic_vector( 16-1 downto 0 );
    a_b_6 : out std_logic_vector( 16-1 downto 0 );
    a_b_7 : out std_logic_vector( 16-1 downto 0 );
    a_b_8 : out std_logic_vector( 16-1 downto 0 );
    a_b_9 : out std_logic_vector( 16-1 downto 0 );
    a_b_10 : out std_logic_vector( 16-1 downto 0 );
    a_b_11 : out std_logic_vector( 16-1 downto 0 );
    a_b_12 : out std_logic_vector( 16-1 downto 0 );
    a_b_13 : out std_logic_vector( 16-1 downto 0 );
    a_b_14 : out std_logic_vector( 16-1 downto 0 );
    a_b_15 : out std_logic_vector( 16-1 downto 0 );
    a_b_16 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_vector_addsub_fabric3;
architecture structural of psb3_0_vector_addsub_fabric3 is 
  signal addsub0_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub3_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub5_s_net : std_logic_vector( 16-1 downto 0 );
  signal mult1_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mult14_p_net : std_logic_vector( 16-1 downto 0 );
  signal addsub8_s_net : std_logic_vector( 16-1 downto 0 );
  signal mult8_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult10_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mult13_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub12_s_net : std_logic_vector( 16-1 downto 0 );
  signal mult0_p_net : std_logic_vector( 16-1 downto 0 );
  signal addsub7_s_net : std_logic_vector( 16-1 downto 0 );
  signal mult6_p_net : std_logic_vector( 16-1 downto 0 );
  signal addsub10_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub14_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub6_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub9_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub13_s_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mult3_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult5_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult7_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult11_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult12_p_net : std_logic_vector( 16-1 downto 0 );
  signal addsub11_s_net : std_logic_vector( 16-1 downto 0 );
  signal mult2_p_net : std_logic_vector( 16-1 downto 0 );
  signal addsub15_s_net : std_logic_vector( 16-1 downto 0 );
  signal mult9_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult15_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult4_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal clk_net : std_logic;
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal ce_net : std_logic;
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
begin
  a_b_1 <= addsub0_s_net;
  a_b_2 <= addsub1_s_net;
  a_b_3 <= addsub2_s_net;
  a_b_4 <= addsub3_s_net;
  a_b_5 <= addsub4_s_net;
  a_b_6 <= addsub5_s_net;
  a_b_7 <= addsub6_s_net;
  a_b_8 <= addsub7_s_net;
  a_b_9 <= addsub8_s_net;
  a_b_10 <= addsub9_s_net;
  a_b_11 <= addsub10_s_net;
  a_b_12 <= addsub11_s_net;
  a_b_13 <= addsub12_s_net;
  a_b_14 <= addsub13_s_net;
  a_b_15 <= addsub14_s_net;
  a_b_16 <= addsub15_s_net;
  mult0_p_net <= a_1;
  reinterpret0_output_port_net <= b_1;
  mult1_p_net <= a_2;
  mult2_p_net <= a_3;
  mult3_p_net <= a_4;
  mult4_p_net <= a_5;
  mult5_p_net <= a_6;
  mult6_p_net <= a_7;
  mult7_p_net <= a_8;
  mult8_p_net <= a_9;
  mult9_p_net <= a_10;
  mult10_p_net <= a_11;
  mult11_p_net <= a_12;
  mult12_p_net <= a_13;
  mult13_p_net <= a_14;
  mult14_p_net <= a_15;
  mult15_p_net <= a_16;
  reinterpret1_output_port_net <= b_2;
  reinterpret2_output_port_net <= b_3;
  reinterpret3_output_port_net <= b_4;
  reinterpret4_output_port_net <= b_5;
  reinterpret5_output_port_net <= b_6;
  reinterpret6_output_port_net <= b_7;
  reinterpret7_output_port_net <= b_8;
  reinterpret8_output_port_net <= b_9;
  reinterpret9_output_port_net <= b_10;
  reinterpret10_output_port_net <= b_11;
  reinterpret11_output_port_net <= b_12;
  reinterpret12_output_port_net <= b_13;
  reinterpret13_output_port_net <= b_14;
  reinterpret14_output_port_net <= b_15;
  reinterpret15_output_port_net <= b_16;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub0 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult0_p_net,
    b => reinterpret0_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub0_s_net
  );
  addsub1 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult1_p_net,
    b => reinterpret1_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  addsub2 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult2_p_net,
    b => reinterpret2_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub2_s_net
  );
  addsub3 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult3_p_net,
    b => reinterpret3_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub3_s_net
  );
  addsub4 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult4_p_net,
    b => reinterpret4_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub4_s_net
  );
  addsub5 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult5_p_net,
    b => reinterpret5_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub5_s_net
  );
  addsub6 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult6_p_net,
    b => reinterpret6_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub6_s_net
  );
  addsub7 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult7_p_net,
    b => reinterpret7_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub7_s_net
  );
  addsub8 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult8_p_net,
    b => reinterpret8_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub8_s_net
  );
  addsub9 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult9_p_net,
    b => reinterpret9_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub9_s_net
  );
  addsub10 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult10_p_net,
    b => reinterpret10_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub10_s_net
  );
  addsub11 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult11_p_net,
    b => reinterpret11_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub11_s_net
  );
  addsub12 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult12_p_net,
    b => reinterpret12_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub12_s_net
  );
  addsub13 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult13_p_net,
    b => reinterpret13_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub13_s_net
  );
  addsub14 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult14_p_net,
    b => reinterpret14_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub14_s_net
  );
  addsub15 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult15_p_net,
    b => reinterpret15_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub15_s_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Vector AddSub Fabric4
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_addsub_fabric4 is
  port (
    a_1 : in std_logic_vector( 16-1 downto 0 );
    b_1 : in std_logic_vector( 16-1 downto 0 );
    a_2 : in std_logic_vector( 16-1 downto 0 );
    a_3 : in std_logic_vector( 16-1 downto 0 );
    a_4 : in std_logic_vector( 16-1 downto 0 );
    a_5 : in std_logic_vector( 16-1 downto 0 );
    a_6 : in std_logic_vector( 16-1 downto 0 );
    a_7 : in std_logic_vector( 16-1 downto 0 );
    a_8 : in std_logic_vector( 16-1 downto 0 );
    a_9 : in std_logic_vector( 16-1 downto 0 );
    a_10 : in std_logic_vector( 16-1 downto 0 );
    a_11 : in std_logic_vector( 16-1 downto 0 );
    a_12 : in std_logic_vector( 16-1 downto 0 );
    a_13 : in std_logic_vector( 16-1 downto 0 );
    a_14 : in std_logic_vector( 16-1 downto 0 );
    a_15 : in std_logic_vector( 16-1 downto 0 );
    a_16 : in std_logic_vector( 16-1 downto 0 );
    b_2 : in std_logic_vector( 16-1 downto 0 );
    b_3 : in std_logic_vector( 16-1 downto 0 );
    b_4 : in std_logic_vector( 16-1 downto 0 );
    b_5 : in std_logic_vector( 16-1 downto 0 );
    b_6 : in std_logic_vector( 16-1 downto 0 );
    b_7 : in std_logic_vector( 16-1 downto 0 );
    b_8 : in std_logic_vector( 16-1 downto 0 );
    b_9 : in std_logic_vector( 16-1 downto 0 );
    b_10 : in std_logic_vector( 16-1 downto 0 );
    b_11 : in std_logic_vector( 16-1 downto 0 );
    b_12 : in std_logic_vector( 16-1 downto 0 );
    b_13 : in std_logic_vector( 16-1 downto 0 );
    b_14 : in std_logic_vector( 16-1 downto 0 );
    b_15 : in std_logic_vector( 16-1 downto 0 );
    b_16 : in std_logic_vector( 16-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    a_b_1 : out std_logic_vector( 16-1 downto 0 );
    a_b_2 : out std_logic_vector( 16-1 downto 0 );
    a_b_3 : out std_logic_vector( 16-1 downto 0 );
    a_b_4 : out std_logic_vector( 16-1 downto 0 );
    a_b_5 : out std_logic_vector( 16-1 downto 0 );
    a_b_6 : out std_logic_vector( 16-1 downto 0 );
    a_b_7 : out std_logic_vector( 16-1 downto 0 );
    a_b_8 : out std_logic_vector( 16-1 downto 0 );
    a_b_9 : out std_logic_vector( 16-1 downto 0 );
    a_b_10 : out std_logic_vector( 16-1 downto 0 );
    a_b_11 : out std_logic_vector( 16-1 downto 0 );
    a_b_12 : out std_logic_vector( 16-1 downto 0 );
    a_b_13 : out std_logic_vector( 16-1 downto 0 );
    a_b_14 : out std_logic_vector( 16-1 downto 0 );
    a_b_15 : out std_logic_vector( 16-1 downto 0 );
    a_b_16 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_vector_addsub_fabric4;
architecture structural of psb3_0_vector_addsub_fabric4 is 
  signal mult8_p_net : std_logic_vector( 16-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub10_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 16-1 downto 0 );
  signal mult10_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult1_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult9_p_net : std_logic_vector( 16-1 downto 0 );
  signal addsub12_s_net : std_logic_vector( 16-1 downto 0 );
  signal mult0_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult3_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult5_p_net : std_logic_vector( 16-1 downto 0 );
  signal addsub3_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub15_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub6_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub0_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub5_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub11_s_net : std_logic_vector( 16-1 downto 0 );
  signal mult6_p_net : std_logic_vector( 16-1 downto 0 );
  signal addsub9_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub14_s_net : std_logic_vector( 16-1 downto 0 );
  signal mult2_p_net : std_logic_vector( 16-1 downto 0 );
  signal addsub7_s_net : std_logic_vector( 16-1 downto 0 );
  signal mult7_p_net : std_logic_vector( 16-1 downto 0 );
  signal addsub8_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub13_s_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mult4_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mult14_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mult12_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult13_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mult15_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal clk_net : std_logic;
  signal ce_net : std_logic;
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mult11_p_net : std_logic_vector( 16-1 downto 0 );
begin
  a_b_1 <= addsub0_s_net;
  a_b_2 <= addsub1_s_net;
  a_b_3 <= addsub2_s_net;
  a_b_4 <= addsub3_s_net;
  a_b_5 <= addsub4_s_net;
  a_b_6 <= addsub5_s_net;
  a_b_7 <= addsub6_s_net;
  a_b_8 <= addsub7_s_net;
  a_b_9 <= addsub8_s_net;
  a_b_10 <= addsub9_s_net;
  a_b_11 <= addsub10_s_net;
  a_b_12 <= addsub11_s_net;
  a_b_13 <= addsub12_s_net;
  a_b_14 <= addsub13_s_net;
  a_b_15 <= addsub14_s_net;
  a_b_16 <= addsub15_s_net;
  mult0_p_net <= a_1;
  reinterpret0_output_port_net <= b_1;
  mult1_p_net <= a_2;
  mult2_p_net <= a_3;
  mult3_p_net <= a_4;
  mult4_p_net <= a_5;
  mult5_p_net <= a_6;
  mult6_p_net <= a_7;
  mult7_p_net <= a_8;
  mult8_p_net <= a_9;
  mult9_p_net <= a_10;
  mult10_p_net <= a_11;
  mult11_p_net <= a_12;
  mult12_p_net <= a_13;
  mult13_p_net <= a_14;
  mult14_p_net <= a_15;
  mult15_p_net <= a_16;
  reinterpret1_output_port_net <= b_2;
  reinterpret2_output_port_net <= b_3;
  reinterpret3_output_port_net <= b_4;
  reinterpret4_output_port_net <= b_5;
  reinterpret5_output_port_net <= b_6;
  reinterpret6_output_port_net <= b_7;
  reinterpret7_output_port_net <= b_8;
  reinterpret8_output_port_net <= b_9;
  reinterpret9_output_port_net <= b_10;
  reinterpret10_output_port_net <= b_11;
  reinterpret11_output_port_net <= b_12;
  reinterpret12_output_port_net <= b_13;
  reinterpret13_output_port_net <= b_14;
  reinterpret14_output_port_net <= b_15;
  reinterpret15_output_port_net <= b_16;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub0 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult0_p_net,
    b => reinterpret0_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub0_s_net
  );
  addsub1 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult1_p_net,
    b => reinterpret1_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  addsub2 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult2_p_net,
    b => reinterpret2_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub2_s_net
  );
  addsub3 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult3_p_net,
    b => reinterpret3_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub3_s_net
  );
  addsub4 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult4_p_net,
    b => reinterpret4_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub4_s_net
  );
  addsub5 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult5_p_net,
    b => reinterpret5_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub5_s_net
  );
  addsub6 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult6_p_net,
    b => reinterpret6_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub6_s_net
  );
  addsub7 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult7_p_net,
    b => reinterpret7_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub7_s_net
  );
  addsub8 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult8_p_net,
    b => reinterpret8_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub8_s_net
  );
  addsub9 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult9_p_net,
    b => reinterpret9_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub9_s_net
  );
  addsub10 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult10_p_net,
    b => reinterpret10_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub10_s_net
  );
  addsub11 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult11_p_net,
    b => reinterpret11_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub11_s_net
  );
  addsub12 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult12_p_net,
    b => reinterpret12_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub12_s_net
  );
  addsub13 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult13_p_net,
    b => reinterpret13_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub13_s_net
  );
  addsub14 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult14_p_net,
    b => reinterpret14_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub14_s_net
  );
  addsub15 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult15_p_net,
    b => reinterpret15_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub15_s_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Vector AddSub Fabric5
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_addsub_fabric5 is
  port (
    a_1 : in std_logic_vector( 16-1 downto 0 );
    b_1 : in std_logic_vector( 16-1 downto 0 );
    a_2 : in std_logic_vector( 16-1 downto 0 );
    a_3 : in std_logic_vector( 16-1 downto 0 );
    a_4 : in std_logic_vector( 16-1 downto 0 );
    a_5 : in std_logic_vector( 16-1 downto 0 );
    a_6 : in std_logic_vector( 16-1 downto 0 );
    a_7 : in std_logic_vector( 16-1 downto 0 );
    a_8 : in std_logic_vector( 16-1 downto 0 );
    a_9 : in std_logic_vector( 16-1 downto 0 );
    a_10 : in std_logic_vector( 16-1 downto 0 );
    a_11 : in std_logic_vector( 16-1 downto 0 );
    a_12 : in std_logic_vector( 16-1 downto 0 );
    a_13 : in std_logic_vector( 16-1 downto 0 );
    a_14 : in std_logic_vector( 16-1 downto 0 );
    a_15 : in std_logic_vector( 16-1 downto 0 );
    a_16 : in std_logic_vector( 16-1 downto 0 );
    b_2 : in std_logic_vector( 16-1 downto 0 );
    b_3 : in std_logic_vector( 16-1 downto 0 );
    b_4 : in std_logic_vector( 16-1 downto 0 );
    b_5 : in std_logic_vector( 16-1 downto 0 );
    b_6 : in std_logic_vector( 16-1 downto 0 );
    b_7 : in std_logic_vector( 16-1 downto 0 );
    b_8 : in std_logic_vector( 16-1 downto 0 );
    b_9 : in std_logic_vector( 16-1 downto 0 );
    b_10 : in std_logic_vector( 16-1 downto 0 );
    b_11 : in std_logic_vector( 16-1 downto 0 );
    b_12 : in std_logic_vector( 16-1 downto 0 );
    b_13 : in std_logic_vector( 16-1 downto 0 );
    b_14 : in std_logic_vector( 16-1 downto 0 );
    b_15 : in std_logic_vector( 16-1 downto 0 );
    b_16 : in std_logic_vector( 16-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    a_b_1 : out std_logic_vector( 16-1 downto 0 );
    a_b_2 : out std_logic_vector( 16-1 downto 0 );
    a_b_3 : out std_logic_vector( 16-1 downto 0 );
    a_b_4 : out std_logic_vector( 16-1 downto 0 );
    a_b_5 : out std_logic_vector( 16-1 downto 0 );
    a_b_6 : out std_logic_vector( 16-1 downto 0 );
    a_b_7 : out std_logic_vector( 16-1 downto 0 );
    a_b_8 : out std_logic_vector( 16-1 downto 0 );
    a_b_9 : out std_logic_vector( 16-1 downto 0 );
    a_b_10 : out std_logic_vector( 16-1 downto 0 );
    a_b_11 : out std_logic_vector( 16-1 downto 0 );
    a_b_12 : out std_logic_vector( 16-1 downto 0 );
    a_b_13 : out std_logic_vector( 16-1 downto 0 );
    a_b_14 : out std_logic_vector( 16-1 downto 0 );
    a_b_15 : out std_logic_vector( 16-1 downto 0 );
    a_b_16 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_vector_addsub_fabric5;
architecture structural of psb3_0_vector_addsub_fabric5 is 
  signal addsub12_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub13_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub14_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub15_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub3_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub5_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub6_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub7_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub0_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub8_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub9_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub11_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub10_s_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mult15_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult10_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult12_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mult4_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult6_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult3_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult9_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mult1_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mult8_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mult5_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult7_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult0_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mult14_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mult2_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult11_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult13_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal ce_net : std_logic;
  signal clk_net : std_logic;
begin
  a_b_1 <= addsub0_s_net;
  a_b_2 <= addsub1_s_net;
  a_b_3 <= addsub2_s_net;
  a_b_4 <= addsub3_s_net;
  a_b_5 <= addsub4_s_net;
  a_b_6 <= addsub5_s_net;
  a_b_7 <= addsub6_s_net;
  a_b_8 <= addsub7_s_net;
  a_b_9 <= addsub8_s_net;
  a_b_10 <= addsub9_s_net;
  a_b_11 <= addsub10_s_net;
  a_b_12 <= addsub11_s_net;
  a_b_13 <= addsub12_s_net;
  a_b_14 <= addsub13_s_net;
  a_b_15 <= addsub14_s_net;
  a_b_16 <= addsub15_s_net;
  mult0_p_net <= a_1;
  reinterpret0_output_port_net <= b_1;
  mult1_p_net <= a_2;
  mult2_p_net <= a_3;
  mult3_p_net <= a_4;
  mult4_p_net <= a_5;
  mult5_p_net <= a_6;
  mult6_p_net <= a_7;
  mult7_p_net <= a_8;
  mult8_p_net <= a_9;
  mult9_p_net <= a_10;
  mult10_p_net <= a_11;
  mult11_p_net <= a_12;
  mult12_p_net <= a_13;
  mult13_p_net <= a_14;
  mult14_p_net <= a_15;
  mult15_p_net <= a_16;
  reinterpret1_output_port_net <= b_2;
  reinterpret2_output_port_net <= b_3;
  reinterpret3_output_port_net <= b_4;
  reinterpret4_output_port_net <= b_5;
  reinterpret5_output_port_net <= b_6;
  reinterpret6_output_port_net <= b_7;
  reinterpret7_output_port_net <= b_8;
  reinterpret8_output_port_net <= b_9;
  reinterpret9_output_port_net <= b_10;
  reinterpret10_output_port_net <= b_11;
  reinterpret11_output_port_net <= b_12;
  reinterpret12_output_port_net <= b_13;
  reinterpret13_output_port_net <= b_14;
  reinterpret14_output_port_net <= b_15;
  reinterpret15_output_port_net <= b_16;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub0 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult0_p_net,
    b => reinterpret0_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub0_s_net
  );
  addsub1 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult1_p_net,
    b => reinterpret1_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  addsub2 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult2_p_net,
    b => reinterpret2_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub2_s_net
  );
  addsub3 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult3_p_net,
    b => reinterpret3_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub3_s_net
  );
  addsub4 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult4_p_net,
    b => reinterpret4_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub4_s_net
  );
  addsub5 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult5_p_net,
    b => reinterpret5_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub5_s_net
  );
  addsub6 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult6_p_net,
    b => reinterpret6_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub6_s_net
  );
  addsub7 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult7_p_net,
    b => reinterpret7_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub7_s_net
  );
  addsub8 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult8_p_net,
    b => reinterpret8_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub8_s_net
  );
  addsub9 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult9_p_net,
    b => reinterpret9_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub9_s_net
  );
  addsub10 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult10_p_net,
    b => reinterpret10_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub10_s_net
  );
  addsub11 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult11_p_net,
    b => reinterpret11_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub11_s_net
  );
  addsub12 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult12_p_net,
    b => reinterpret12_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub12_s_net
  );
  addsub13 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult13_p_net,
    b => reinterpret13_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub13_s_net
  );
  addsub14 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult14_p_net,
    b => reinterpret14_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub14_s_net
  );
  addsub15 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult15_p_net,
    b => reinterpret15_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub15_s_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Vector AddSub Fabric6
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_addsub_fabric6 is
  port (
    a_1 : in std_logic_vector( 16-1 downto 0 );
    b_1 : in std_logic_vector( 16-1 downto 0 );
    a_2 : in std_logic_vector( 16-1 downto 0 );
    a_3 : in std_logic_vector( 16-1 downto 0 );
    a_4 : in std_logic_vector( 16-1 downto 0 );
    a_5 : in std_logic_vector( 16-1 downto 0 );
    a_6 : in std_logic_vector( 16-1 downto 0 );
    a_7 : in std_logic_vector( 16-1 downto 0 );
    a_8 : in std_logic_vector( 16-1 downto 0 );
    a_9 : in std_logic_vector( 16-1 downto 0 );
    a_10 : in std_logic_vector( 16-1 downto 0 );
    a_11 : in std_logic_vector( 16-1 downto 0 );
    a_12 : in std_logic_vector( 16-1 downto 0 );
    a_13 : in std_logic_vector( 16-1 downto 0 );
    a_14 : in std_logic_vector( 16-1 downto 0 );
    a_15 : in std_logic_vector( 16-1 downto 0 );
    a_16 : in std_logic_vector( 16-1 downto 0 );
    b_2 : in std_logic_vector( 16-1 downto 0 );
    b_3 : in std_logic_vector( 16-1 downto 0 );
    b_4 : in std_logic_vector( 16-1 downto 0 );
    b_5 : in std_logic_vector( 16-1 downto 0 );
    b_6 : in std_logic_vector( 16-1 downto 0 );
    b_7 : in std_logic_vector( 16-1 downto 0 );
    b_8 : in std_logic_vector( 16-1 downto 0 );
    b_9 : in std_logic_vector( 16-1 downto 0 );
    b_10 : in std_logic_vector( 16-1 downto 0 );
    b_11 : in std_logic_vector( 16-1 downto 0 );
    b_12 : in std_logic_vector( 16-1 downto 0 );
    b_13 : in std_logic_vector( 16-1 downto 0 );
    b_14 : in std_logic_vector( 16-1 downto 0 );
    b_15 : in std_logic_vector( 16-1 downto 0 );
    b_16 : in std_logic_vector( 16-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    a_b_1 : out std_logic_vector( 16-1 downto 0 );
    a_b_2 : out std_logic_vector( 16-1 downto 0 );
    a_b_3 : out std_logic_vector( 16-1 downto 0 );
    a_b_4 : out std_logic_vector( 16-1 downto 0 );
    a_b_5 : out std_logic_vector( 16-1 downto 0 );
    a_b_6 : out std_logic_vector( 16-1 downto 0 );
    a_b_7 : out std_logic_vector( 16-1 downto 0 );
    a_b_8 : out std_logic_vector( 16-1 downto 0 );
    a_b_9 : out std_logic_vector( 16-1 downto 0 );
    a_b_10 : out std_logic_vector( 16-1 downto 0 );
    a_b_11 : out std_logic_vector( 16-1 downto 0 );
    a_b_12 : out std_logic_vector( 16-1 downto 0 );
    a_b_13 : out std_logic_vector( 16-1 downto 0 );
    a_b_14 : out std_logic_vector( 16-1 downto 0 );
    a_b_15 : out std_logic_vector( 16-1 downto 0 );
    a_b_16 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_vector_addsub_fabric6;
architecture structural of psb3_0_vector_addsub_fabric6 is 
  signal addsub3_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub5_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub0_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 16-1 downto 0 );
  signal mult7_p_net : std_logic_vector( 16-1 downto 0 );
  signal addsub8_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub13_s_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub9_s_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub15_s_net : std_logic_vector( 16-1 downto 0 );
  signal mult4_p_net : std_logic_vector( 16-1 downto 0 );
  signal addsub6_s_net : std_logic_vector( 16-1 downto 0 );
  signal mult2_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult13_p_net : std_logic_vector( 16-1 downto 0 );
  signal addsub7_s_net : std_logic_vector( 16-1 downto 0 );
  signal mult10_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult0_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult5_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult9_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult1_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult15_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult6_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult12_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult11_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult14_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub14_s_net : std_logic_vector( 16-1 downto 0 );
  signal mult3_p_net : std_logic_vector( 16-1 downto 0 );
  signal addsub12_s_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mult8_p_net : std_logic_vector( 16-1 downto 0 );
  signal addsub10_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub11_s_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal clk_net : std_logic;
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal ce_net : std_logic;
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
begin
  a_b_1 <= addsub0_s_net;
  a_b_2 <= addsub1_s_net;
  a_b_3 <= addsub2_s_net;
  a_b_4 <= addsub3_s_net;
  a_b_5 <= addsub4_s_net;
  a_b_6 <= addsub5_s_net;
  a_b_7 <= addsub6_s_net;
  a_b_8 <= addsub7_s_net;
  a_b_9 <= addsub8_s_net;
  a_b_10 <= addsub9_s_net;
  a_b_11 <= addsub10_s_net;
  a_b_12 <= addsub11_s_net;
  a_b_13 <= addsub12_s_net;
  a_b_14 <= addsub13_s_net;
  a_b_15 <= addsub14_s_net;
  a_b_16 <= addsub15_s_net;
  mult0_p_net <= a_1;
  reinterpret0_output_port_net <= b_1;
  mult1_p_net <= a_2;
  mult2_p_net <= a_3;
  mult3_p_net <= a_4;
  mult4_p_net <= a_5;
  mult5_p_net <= a_6;
  mult6_p_net <= a_7;
  mult7_p_net <= a_8;
  mult8_p_net <= a_9;
  mult9_p_net <= a_10;
  mult10_p_net <= a_11;
  mult11_p_net <= a_12;
  mult12_p_net <= a_13;
  mult13_p_net <= a_14;
  mult14_p_net <= a_15;
  mult15_p_net <= a_16;
  reinterpret1_output_port_net <= b_2;
  reinterpret2_output_port_net <= b_3;
  reinterpret3_output_port_net <= b_4;
  reinterpret4_output_port_net <= b_5;
  reinterpret5_output_port_net <= b_6;
  reinterpret6_output_port_net <= b_7;
  reinterpret7_output_port_net <= b_8;
  reinterpret8_output_port_net <= b_9;
  reinterpret9_output_port_net <= b_10;
  reinterpret10_output_port_net <= b_11;
  reinterpret11_output_port_net <= b_12;
  reinterpret12_output_port_net <= b_13;
  reinterpret13_output_port_net <= b_14;
  reinterpret14_output_port_net <= b_15;
  reinterpret15_output_port_net <= b_16;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub0 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult0_p_net,
    b => reinterpret0_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub0_s_net
  );
  addsub1 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult1_p_net,
    b => reinterpret1_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  addsub2 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult2_p_net,
    b => reinterpret2_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub2_s_net
  );
  addsub3 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult3_p_net,
    b => reinterpret3_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub3_s_net
  );
  addsub4 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult4_p_net,
    b => reinterpret4_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub4_s_net
  );
  addsub5 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult5_p_net,
    b => reinterpret5_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub5_s_net
  );
  addsub6 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult6_p_net,
    b => reinterpret6_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub6_s_net
  );
  addsub7 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult7_p_net,
    b => reinterpret7_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub7_s_net
  );
  addsub8 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult8_p_net,
    b => reinterpret8_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub8_s_net
  );
  addsub9 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult9_p_net,
    b => reinterpret9_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub9_s_net
  );
  addsub10 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult10_p_net,
    b => reinterpret10_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub10_s_net
  );
  addsub11 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult11_p_net,
    b => reinterpret11_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub11_s_net
  );
  addsub12 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult12_p_net,
    b => reinterpret12_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub12_s_net
  );
  addsub13 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult13_p_net,
    b => reinterpret13_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub13_s_net
  );
  addsub14 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult14_p_net,
    b => reinterpret14_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub14_s_net
  );
  addsub15 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult15_p_net,
    b => reinterpret15_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub15_s_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Vector AddSub Fabric7
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_addsub_fabric7 is
  port (
    a_1 : in std_logic_vector( 16-1 downto 0 );
    b_1 : in std_logic_vector( 16-1 downto 0 );
    a_2 : in std_logic_vector( 16-1 downto 0 );
    a_3 : in std_logic_vector( 16-1 downto 0 );
    a_4 : in std_logic_vector( 16-1 downto 0 );
    a_5 : in std_logic_vector( 16-1 downto 0 );
    a_6 : in std_logic_vector( 16-1 downto 0 );
    a_7 : in std_logic_vector( 16-1 downto 0 );
    a_8 : in std_logic_vector( 16-1 downto 0 );
    a_9 : in std_logic_vector( 16-1 downto 0 );
    a_10 : in std_logic_vector( 16-1 downto 0 );
    a_11 : in std_logic_vector( 16-1 downto 0 );
    a_12 : in std_logic_vector( 16-1 downto 0 );
    a_13 : in std_logic_vector( 16-1 downto 0 );
    a_14 : in std_logic_vector( 16-1 downto 0 );
    a_15 : in std_logic_vector( 16-1 downto 0 );
    a_16 : in std_logic_vector( 16-1 downto 0 );
    b_2 : in std_logic_vector( 16-1 downto 0 );
    b_3 : in std_logic_vector( 16-1 downto 0 );
    b_4 : in std_logic_vector( 16-1 downto 0 );
    b_5 : in std_logic_vector( 16-1 downto 0 );
    b_6 : in std_logic_vector( 16-1 downto 0 );
    b_7 : in std_logic_vector( 16-1 downto 0 );
    b_8 : in std_logic_vector( 16-1 downto 0 );
    b_9 : in std_logic_vector( 16-1 downto 0 );
    b_10 : in std_logic_vector( 16-1 downto 0 );
    b_11 : in std_logic_vector( 16-1 downto 0 );
    b_12 : in std_logic_vector( 16-1 downto 0 );
    b_13 : in std_logic_vector( 16-1 downto 0 );
    b_14 : in std_logic_vector( 16-1 downto 0 );
    b_15 : in std_logic_vector( 16-1 downto 0 );
    b_16 : in std_logic_vector( 16-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    a_b_1 : out std_logic_vector( 16-1 downto 0 );
    a_b_2 : out std_logic_vector( 16-1 downto 0 );
    a_b_3 : out std_logic_vector( 16-1 downto 0 );
    a_b_4 : out std_logic_vector( 16-1 downto 0 );
    a_b_5 : out std_logic_vector( 16-1 downto 0 );
    a_b_6 : out std_logic_vector( 16-1 downto 0 );
    a_b_7 : out std_logic_vector( 16-1 downto 0 );
    a_b_8 : out std_logic_vector( 16-1 downto 0 );
    a_b_9 : out std_logic_vector( 16-1 downto 0 );
    a_b_10 : out std_logic_vector( 16-1 downto 0 );
    a_b_11 : out std_logic_vector( 16-1 downto 0 );
    a_b_12 : out std_logic_vector( 16-1 downto 0 );
    a_b_13 : out std_logic_vector( 16-1 downto 0 );
    a_b_14 : out std_logic_vector( 16-1 downto 0 );
    a_b_15 : out std_logic_vector( 16-1 downto 0 );
    a_b_16 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_vector_addsub_fabric7;
architecture structural of psb3_0_vector_addsub_fabric7 is 
  signal addsub10_s_net : std_logic_vector( 16-1 downto 0 );
  signal mult6_p_net : std_logic_vector( 16-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub11_s_net : std_logic_vector( 16-1 downto 0 );
  signal mult7_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult9_p_net : std_logic_vector( 16-1 downto 0 );
  signal addsub15_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub7_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub13_s_net : std_logic_vector( 16-1 downto 0 );
  signal mult0_p_net : std_logic_vector( 16-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 16-1 downto 0 );
  signal mult3_p_net : std_logic_vector( 16-1 downto 0 );
  signal addsub9_s_net : std_logic_vector( 16-1 downto 0 );
  signal mult1_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult5_p_net : std_logic_vector( 16-1 downto 0 );
  signal addsub0_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub6_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub12_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub14_s_net : std_logic_vector( 16-1 downto 0 );
  signal mult8_p_net : std_logic_vector( 16-1 downto 0 );
  signal addsub3_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub8_s_net : std_logic_vector( 16-1 downto 0 );
  signal mult2_p_net : std_logic_vector( 16-1 downto 0 );
  signal addsub5_s_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mult4_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal clk_net : std_logic;
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mult11_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mult13_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal ce_net : std_logic;
  signal mult15_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult12_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult14_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult10_p_net : std_logic_vector( 16-1 downto 0 );
begin
  a_b_1 <= addsub0_s_net;
  a_b_2 <= addsub1_s_net;
  a_b_3 <= addsub2_s_net;
  a_b_4 <= addsub3_s_net;
  a_b_5 <= addsub4_s_net;
  a_b_6 <= addsub5_s_net;
  a_b_7 <= addsub6_s_net;
  a_b_8 <= addsub7_s_net;
  a_b_9 <= addsub8_s_net;
  a_b_10 <= addsub9_s_net;
  a_b_11 <= addsub10_s_net;
  a_b_12 <= addsub11_s_net;
  a_b_13 <= addsub12_s_net;
  a_b_14 <= addsub13_s_net;
  a_b_15 <= addsub14_s_net;
  a_b_16 <= addsub15_s_net;
  mult0_p_net <= a_1;
  reinterpret0_output_port_net <= b_1;
  mult1_p_net <= a_2;
  mult2_p_net <= a_3;
  mult3_p_net <= a_4;
  mult4_p_net <= a_5;
  mult5_p_net <= a_6;
  mult6_p_net <= a_7;
  mult7_p_net <= a_8;
  mult8_p_net <= a_9;
  mult9_p_net <= a_10;
  mult10_p_net <= a_11;
  mult11_p_net <= a_12;
  mult12_p_net <= a_13;
  mult13_p_net <= a_14;
  mult14_p_net <= a_15;
  mult15_p_net <= a_16;
  reinterpret1_output_port_net <= b_2;
  reinterpret2_output_port_net <= b_3;
  reinterpret3_output_port_net <= b_4;
  reinterpret4_output_port_net <= b_5;
  reinterpret5_output_port_net <= b_6;
  reinterpret6_output_port_net <= b_7;
  reinterpret7_output_port_net <= b_8;
  reinterpret8_output_port_net <= b_9;
  reinterpret9_output_port_net <= b_10;
  reinterpret10_output_port_net <= b_11;
  reinterpret11_output_port_net <= b_12;
  reinterpret12_output_port_net <= b_13;
  reinterpret13_output_port_net <= b_14;
  reinterpret14_output_port_net <= b_15;
  reinterpret15_output_port_net <= b_16;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub0 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult0_p_net,
    b => reinterpret0_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub0_s_net
  );
  addsub1 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult1_p_net,
    b => reinterpret1_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  addsub2 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult2_p_net,
    b => reinterpret2_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub2_s_net
  );
  addsub3 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult3_p_net,
    b => reinterpret3_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub3_s_net
  );
  addsub4 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult4_p_net,
    b => reinterpret4_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub4_s_net
  );
  addsub5 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult5_p_net,
    b => reinterpret5_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub5_s_net
  );
  addsub6 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult6_p_net,
    b => reinterpret6_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub6_s_net
  );
  addsub7 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult7_p_net,
    b => reinterpret7_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub7_s_net
  );
  addsub8 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult8_p_net,
    b => reinterpret8_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub8_s_net
  );
  addsub9 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult9_p_net,
    b => reinterpret9_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub9_s_net
  );
  addsub10 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult10_p_net,
    b => reinterpret10_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub10_s_net
  );
  addsub11 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult11_p_net,
    b => reinterpret11_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub11_s_net
  );
  addsub12 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult12_p_net,
    b => reinterpret12_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub12_s_net
  );
  addsub13 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult13_p_net,
    b => reinterpret13_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub13_s_net
  );
  addsub14 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult14_p_net,
    b => reinterpret14_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub14_s_net
  );
  addsub15 : entity xil_defaultlib.psb3_0_xladdsub 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 14,
    b_width => 16,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 18,
    core_name0 => "psb3_0_c_addsub_v12_0_i2",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 18,
    latency => 2,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 14,
    s_width => 16
  )
  port map (
    clr => '0',
    en => "1",
    a => mult15_p_net,
    b => reinterpret15_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub15_s_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Vector Constant
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_constant is
  port (
    out1_1 : out std_logic_vector( 16-1 downto 0 );
    out1_2 : out std_logic_vector( 16-1 downto 0 );
    out1_3 : out std_logic_vector( 16-1 downto 0 );
    out1_4 : out std_logic_vector( 16-1 downto 0 );
    out1_5 : out std_logic_vector( 16-1 downto 0 );
    out1_6 : out std_logic_vector( 16-1 downto 0 );
    out1_7 : out std_logic_vector( 16-1 downto 0 );
    out1_8 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_vector_constant;
architecture structural of psb3_0_vector_constant is 
  signal constant7_op_net : std_logic_vector( 16-1 downto 0 );
  signal constant3_op_net : std_logic_vector( 16-1 downto 0 );
  signal constant6_op_net : std_logic_vector( 16-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 16-1 downto 0 );
  signal constant2_op_net : std_logic_vector( 16-1 downto 0 );
  signal constant5_op_net : std_logic_vector( 16-1 downto 0 );
  signal constant4_op_net : std_logic_vector( 16-1 downto 0 );
  signal constant0_op_net : std_logic_vector( 16-1 downto 0 );
begin
  out1_1 <= constant0_op_net;
  out1_2 <= constant1_op_net;
  out1_3 <= constant2_op_net;
  out1_4 <= constant3_op_net;
  out1_5 <= constant4_op_net;
  out1_6 <= constant5_op_net;
  out1_7 <= constant6_op_net;
  out1_8 <= constant7_op_net;
  constant0 : entity xil_defaultlib.sysgen_constant_53872fb2be 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant0_op_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_53872fb2be 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  constant2 : entity xil_defaultlib.sysgen_constant_53872fb2be 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant2_op_net
  );
  constant3 : entity xil_defaultlib.sysgen_constant_53872fb2be 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant3_op_net
  );
  constant4 : entity xil_defaultlib.sysgen_constant_53872fb2be 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant4_op_net
  );
  constant5 : entity xil_defaultlib.sysgen_constant_53872fb2be 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant5_op_net
  );
  constant6 : entity xil_defaultlib.sysgen_constant_53872fb2be 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant6_op_net
  );
  constant7 : entity xil_defaultlib.sysgen_constant_53872fb2be 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant7_op_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Vector Mux
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_mux is
  port (
    sel : in std_logic_vector( 1-1 downto 0 );
    i0_1 : in std_logic_vector( 16-1 downto 0 );
    i1_1 : in std_logic_vector( 20-1 downto 0 );
    i0_2 : in std_logic_vector( 16-1 downto 0 );
    i0_3 : in std_logic_vector( 16-1 downto 0 );
    i0_4 : in std_logic_vector( 16-1 downto 0 );
    i0_5 : in std_logic_vector( 16-1 downto 0 );
    i0_6 : in std_logic_vector( 16-1 downto 0 );
    i0_7 : in std_logic_vector( 16-1 downto 0 );
    i0_8 : in std_logic_vector( 16-1 downto 0 );
    i1_2 : in std_logic_vector( 20-1 downto 0 );
    i1_3 : in std_logic_vector( 20-1 downto 0 );
    i1_4 : in std_logic_vector( 20-1 downto 0 );
    i1_5 : in std_logic_vector( 20-1 downto 0 );
    i1_6 : in std_logic_vector( 20-1 downto 0 );
    i1_7 : in std_logic_vector( 20-1 downto 0 );
    i1_8 : in std_logic_vector( 20-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    o_1 : out std_logic_vector( 16-1 downto 0 );
    o_2 : out std_logic_vector( 16-1 downto 0 );
    o_3 : out std_logic_vector( 16-1 downto 0 );
    o_4 : out std_logic_vector( 16-1 downto 0 );
    o_5 : out std_logic_vector( 16-1 downto 0 );
    o_6 : out std_logic_vector( 16-1 downto 0 );
    o_7 : out std_logic_vector( 16-1 downto 0 );
    o_8 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_vector_mux;
architecture structural of psb3_0_vector_mux is 
  signal reinterpret27_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 16-1 downto 0 );
  signal mux6_y_net : std_logic_vector( 16-1 downto 0 );
  signal constant2_op_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret29_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal reinterpret24_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret30_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal mux2_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret25_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal constant7_op_net : std_logic_vector( 16-1 downto 0 );
  signal mux4_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret26_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal register_q_net : std_logic_vector( 1-1 downto 0 );
  signal constant5_op_net : std_logic_vector( 16-1 downto 0 );
  signal mux0_y_net : std_logic_vector( 16-1 downto 0 );
  signal mux5_y_net : std_logic_vector( 16-1 downto 0 );
  signal mux3_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret28_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal constant3_op_net : std_logic_vector( 16-1 downto 0 );
  signal constant4_op_net : std_logic_vector( 16-1 downto 0 );
  signal constant0_op_net : std_logic_vector( 16-1 downto 0 );
  signal mux7_y_net : std_logic_vector( 16-1 downto 0 );
  signal constant6_op_net : std_logic_vector( 16-1 downto 0 );
  signal ce_net : std_logic;
  signal reinterpret31_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal clk_net : std_logic;
begin
  o_1 <= mux0_y_net;
  o_2 <= mux1_y_net;
  o_3 <= mux2_y_net;
  o_4 <= mux3_y_net;
  o_5 <= mux4_y_net;
  o_6 <= mux5_y_net;
  o_7 <= mux6_y_net;
  o_8 <= mux7_y_net;
  register_q_net <= sel;
  constant0_op_net <= i0_1;
  reinterpret24_output_port_net <= i1_1;
  constant1_op_net <= i0_2;
  constant2_op_net <= i0_3;
  constant3_op_net <= i0_4;
  constant4_op_net <= i0_5;
  constant5_op_net <= i0_6;
  constant6_op_net <= i0_7;
  constant7_op_net <= i0_8;
  reinterpret25_output_port_net <= i1_2;
  reinterpret26_output_port_net <= i1_3;
  reinterpret27_output_port_net <= i1_4;
  reinterpret28_output_port_net <= i1_5;
  reinterpret29_output_port_net <= i1_6;
  reinterpret30_output_port_net <= i1_7;
  reinterpret31_output_port_net <= i1_8;
  clk_net <= clk_1;
  ce_net <= ce_1;
  mux0 : entity xil_defaultlib.sysgen_mux_7ec6aa7932 
  port map (
    clr => '0',
    sel => register_q_net,
    d0 => constant0_op_net,
    d1 => reinterpret24_output_port_net,
    clk => clk_net,
    ce => ce_net,
    y => mux0_y_net
  );
  mux1 : entity xil_defaultlib.sysgen_mux_7ec6aa7932 
  port map (
    clr => '0',
    sel => register_q_net,
    d0 => constant1_op_net,
    d1 => reinterpret25_output_port_net,
    clk => clk_net,
    ce => ce_net,
    y => mux1_y_net
  );
  mux2 : entity xil_defaultlib.sysgen_mux_7ec6aa7932 
  port map (
    clr => '0',
    sel => register_q_net,
    d0 => constant2_op_net,
    d1 => reinterpret26_output_port_net,
    clk => clk_net,
    ce => ce_net,
    y => mux2_y_net
  );
  mux3 : entity xil_defaultlib.sysgen_mux_7ec6aa7932 
  port map (
    clr => '0',
    sel => register_q_net,
    d0 => constant3_op_net,
    d1 => reinterpret27_output_port_net,
    clk => clk_net,
    ce => ce_net,
    y => mux3_y_net
  );
  mux4 : entity xil_defaultlib.sysgen_mux_7ec6aa7932 
  port map (
    clr => '0',
    sel => register_q_net,
    d0 => constant4_op_net,
    d1 => reinterpret28_output_port_net,
    clk => clk_net,
    ce => ce_net,
    y => mux4_y_net
  );
  mux5 : entity xil_defaultlib.sysgen_mux_7ec6aa7932 
  port map (
    clr => '0',
    sel => register_q_net,
    d0 => constant5_op_net,
    d1 => reinterpret29_output_port_net,
    clk => clk_net,
    ce => ce_net,
    y => mux5_y_net
  );
  mux6 : entity xil_defaultlib.sysgen_mux_7ec6aa7932 
  port map (
    clr => '0',
    sel => register_q_net,
    d0 => constant6_op_net,
    d1 => reinterpret30_output_port_net,
    clk => clk_net,
    ce => ce_net,
    y => mux6_y_net
  );
  mux7 : entity xil_defaultlib.sysgen_mux_7ec6aa7932 
  port map (
    clr => '0',
    sel => register_q_net,
    d0 => constant7_op_net,
    d1 => reinterpret31_output_port_net,
    clk => clk_net,
    ce => ce_net,
    y => mux7_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Vector Mux1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_mux1 is
  port (
    sel : in std_logic_vector( 1-1 downto 0 );
    i0_1 : in std_logic_vector( 16-1 downto 0 );
    i1_1 : in std_logic_vector( 20-1 downto 0 );
    i0_2 : in std_logic_vector( 16-1 downto 0 );
    i0_3 : in std_logic_vector( 16-1 downto 0 );
    i0_4 : in std_logic_vector( 16-1 downto 0 );
    i0_5 : in std_logic_vector( 16-1 downto 0 );
    i0_6 : in std_logic_vector( 16-1 downto 0 );
    i0_7 : in std_logic_vector( 16-1 downto 0 );
    i0_8 : in std_logic_vector( 16-1 downto 0 );
    i1_2 : in std_logic_vector( 20-1 downto 0 );
    i1_3 : in std_logic_vector( 20-1 downto 0 );
    i1_4 : in std_logic_vector( 20-1 downto 0 );
    i1_5 : in std_logic_vector( 20-1 downto 0 );
    i1_6 : in std_logic_vector( 20-1 downto 0 );
    i1_7 : in std_logic_vector( 20-1 downto 0 );
    i1_8 : in std_logic_vector( 20-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    o_1 : out std_logic_vector( 16-1 downto 0 );
    o_2 : out std_logic_vector( 16-1 downto 0 );
    o_3 : out std_logic_vector( 16-1 downto 0 );
    o_4 : out std_logic_vector( 16-1 downto 0 );
    o_5 : out std_logic_vector( 16-1 downto 0 );
    o_6 : out std_logic_vector( 16-1 downto 0 );
    o_7 : out std_logic_vector( 16-1 downto 0 );
    o_8 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_vector_mux1;
architecture structural of psb3_0_vector_mux1 is 
  signal mux0_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret17_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal reinterpret20_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal clk_net : std_logic;
  signal ce_net : std_logic;
  signal constant3_op_net : std_logic_vector( 16-1 downto 0 );
  signal mux6_y_net : std_logic_vector( 16-1 downto 0 );
  signal constant6_op_net : std_logic_vector( 16-1 downto 0 );
  signal constant4_op_net : std_logic_vector( 16-1 downto 0 );
  signal mux3_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret18_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal constant0_op_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret22_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal reinterpret16_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal mux5_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret23_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 16-1 downto 0 );
  signal mux4_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret19_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal mux2_y_net : std_logic_vector( 16-1 downto 0 );
  signal constant5_op_net : std_logic_vector( 16-1 downto 0 );
  signal mux7_y_net : std_logic_vector( 16-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 16-1 downto 0 );
  signal constant7_op_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret21_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal register_q_net : std_logic_vector( 1-1 downto 0 );
  signal constant2_op_net : std_logic_vector( 16-1 downto 0 );
begin
  o_1 <= mux0_y_net;
  o_2 <= mux1_y_net;
  o_3 <= mux2_y_net;
  o_4 <= mux3_y_net;
  o_5 <= mux4_y_net;
  o_6 <= mux5_y_net;
  o_7 <= mux6_y_net;
  o_8 <= mux7_y_net;
  register_q_net <= sel;
  constant0_op_net <= i0_1;
  reinterpret16_output_port_net <= i1_1;
  constant1_op_net <= i0_2;
  constant2_op_net <= i0_3;
  constant3_op_net <= i0_4;
  constant4_op_net <= i0_5;
  constant5_op_net <= i0_6;
  constant6_op_net <= i0_7;
  constant7_op_net <= i0_8;
  reinterpret17_output_port_net <= i1_2;
  reinterpret18_output_port_net <= i1_3;
  reinterpret19_output_port_net <= i1_4;
  reinterpret20_output_port_net <= i1_5;
  reinterpret21_output_port_net <= i1_6;
  reinterpret22_output_port_net <= i1_7;
  reinterpret23_output_port_net <= i1_8;
  clk_net <= clk_1;
  ce_net <= ce_1;
  mux0 : entity xil_defaultlib.sysgen_mux_7ec6aa7932 
  port map (
    clr => '0',
    sel => register_q_net,
    d0 => constant0_op_net,
    d1 => reinterpret16_output_port_net,
    clk => clk_net,
    ce => ce_net,
    y => mux0_y_net
  );
  mux1 : entity xil_defaultlib.sysgen_mux_7ec6aa7932 
  port map (
    clr => '0',
    sel => register_q_net,
    d0 => constant1_op_net,
    d1 => reinterpret17_output_port_net,
    clk => clk_net,
    ce => ce_net,
    y => mux1_y_net
  );
  mux2 : entity xil_defaultlib.sysgen_mux_7ec6aa7932 
  port map (
    clr => '0',
    sel => register_q_net,
    d0 => constant2_op_net,
    d1 => reinterpret18_output_port_net,
    clk => clk_net,
    ce => ce_net,
    y => mux2_y_net
  );
  mux3 : entity xil_defaultlib.sysgen_mux_7ec6aa7932 
  port map (
    clr => '0',
    sel => register_q_net,
    d0 => constant3_op_net,
    d1 => reinterpret19_output_port_net,
    clk => clk_net,
    ce => ce_net,
    y => mux3_y_net
  );
  mux4 : entity xil_defaultlib.sysgen_mux_7ec6aa7932 
  port map (
    clr => '0',
    sel => register_q_net,
    d0 => constant4_op_net,
    d1 => reinterpret20_output_port_net,
    clk => clk_net,
    ce => ce_net,
    y => mux4_y_net
  );
  mux5 : entity xil_defaultlib.sysgen_mux_7ec6aa7932 
  port map (
    clr => '0',
    sel => register_q_net,
    d0 => constant5_op_net,
    d1 => reinterpret21_output_port_net,
    clk => clk_net,
    ce => ce_net,
    y => mux5_y_net
  );
  mux6 : entity xil_defaultlib.sysgen_mux_7ec6aa7932 
  port map (
    clr => '0',
    sel => register_q_net,
    d0 => constant6_op_net,
    d1 => reinterpret22_output_port_net,
    clk => clk_net,
    ce => ce_net,
    y => mux6_y_net
  );
  mux7 : entity xil_defaultlib.sysgen_mux_7ec6aa7932 
  port map (
    clr => '0',
    sel => register_q_net,
    d0 => constant7_op_net,
    d1 => reinterpret23_output_port_net,
    clk => clk_net,
    ce => ce_net,
    y => mux7_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Vector Real Mult Im_1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_real_mult_im_1 is
  port (
    a_1 : in std_logic_vector( 16-1 downto 0 );
    b_1 : in std_logic_vector( 16-1 downto 0 );
    a_2 : in std_logic_vector( 16-1 downto 0 );
    a_3 : in std_logic_vector( 16-1 downto 0 );
    a_4 : in std_logic_vector( 16-1 downto 0 );
    a_5 : in std_logic_vector( 16-1 downto 0 );
    a_6 : in std_logic_vector( 16-1 downto 0 );
    a_7 : in std_logic_vector( 16-1 downto 0 );
    a_8 : in std_logic_vector( 16-1 downto 0 );
    a_9 : in std_logic_vector( 16-1 downto 0 );
    a_10 : in std_logic_vector( 16-1 downto 0 );
    a_11 : in std_logic_vector( 16-1 downto 0 );
    a_12 : in std_logic_vector( 16-1 downto 0 );
    a_13 : in std_logic_vector( 16-1 downto 0 );
    a_14 : in std_logic_vector( 16-1 downto 0 );
    a_15 : in std_logic_vector( 16-1 downto 0 );
    a_16 : in std_logic_vector( 16-1 downto 0 );
    b_2 : in std_logic_vector( 16-1 downto 0 );
    b_3 : in std_logic_vector( 16-1 downto 0 );
    b_4 : in std_logic_vector( 16-1 downto 0 );
    b_5 : in std_logic_vector( 16-1 downto 0 );
    b_6 : in std_logic_vector( 16-1 downto 0 );
    b_7 : in std_logic_vector( 16-1 downto 0 );
    b_8 : in std_logic_vector( 16-1 downto 0 );
    b_9 : in std_logic_vector( 16-1 downto 0 );
    b_10 : in std_logic_vector( 16-1 downto 0 );
    b_11 : in std_logic_vector( 16-1 downto 0 );
    b_12 : in std_logic_vector( 16-1 downto 0 );
    b_13 : in std_logic_vector( 16-1 downto 0 );
    b_14 : in std_logic_vector( 16-1 downto 0 );
    b_15 : in std_logic_vector( 16-1 downto 0 );
    b_16 : in std_logic_vector( 16-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    a_x_b_1 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_2 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_3 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_4 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_5 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_6 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_7 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_8 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_9 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_10 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_11 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_12 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_13 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_14 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_15 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_16 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_vector_real_mult_im_1;
architecture structural of psb3_0_vector_real_mult_im_1 is 
  signal mult5_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult6_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult4_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult7_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult8_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult0_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult1_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult2_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult3_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal mult15_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mult9_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult14_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult11_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mult13_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal mult12_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal mult10_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal clk_net : std_logic;
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal ce_net : std_logic;
begin
  a_x_b_1 <= mult0_p_net;
  a_x_b_2 <= mult1_p_net;
  a_x_b_3 <= mult2_p_net;
  a_x_b_4 <= mult3_p_net;
  a_x_b_5 <= mult4_p_net;
  a_x_b_6 <= mult5_p_net;
  a_x_b_7 <= mult6_p_net;
  a_x_b_8 <= mult7_p_net;
  a_x_b_9 <= mult8_p_net;
  a_x_b_10 <= mult9_p_net;
  a_x_b_11 <= mult10_p_net;
  a_x_b_12 <= mult11_p_net;
  a_x_b_13 <= mult12_p_net;
  a_x_b_14 <= mult13_p_net;
  a_x_b_15 <= mult14_p_net;
  a_x_b_16 <= mult15_p_net;
  reinterpret0_output_port_net <= a_1;
  reinterpret0_output_port_net_x0 <= b_1;
  reinterpret1_output_port_net <= a_2;
  reinterpret2_output_port_net_x0 <= a_3;
  reinterpret3_output_port_net_x0 <= a_4;
  reinterpret4_output_port_net <= a_5;
  reinterpret5_output_port_net_x0 <= a_6;
  reinterpret6_output_port_net <= a_7;
  reinterpret7_output_port_net_x0 <= a_8;
  reinterpret8_output_port_net_x0 <= a_9;
  reinterpret9_output_port_net_x0 <= a_10;
  reinterpret10_output_port_net_x0 <= a_11;
  reinterpret11_output_port_net_x0 <= a_12;
  reinterpret12_output_port_net_x0 <= a_13;
  reinterpret13_output_port_net_x0 <= a_14;
  reinterpret14_output_port_net_x0 <= a_15;
  reinterpret15_output_port_net_x0 <= a_16;
  reinterpret1_output_port_net_x0 <= b_2;
  reinterpret2_output_port_net <= b_3;
  reinterpret3_output_port_net <= b_4;
  reinterpret4_output_port_net_x0 <= b_5;
  reinterpret5_output_port_net <= b_6;
  reinterpret6_output_port_net_x0 <= b_7;
  reinterpret7_output_port_net <= b_8;
  reinterpret8_output_port_net <= b_9;
  reinterpret9_output_port_net <= b_10;
  reinterpret10_output_port_net <= b_11;
  reinterpret11_output_port_net <= b_12;
  reinterpret12_output_port_net <= b_13;
  reinterpret13_output_port_net <= b_14;
  reinterpret14_output_port_net <= b_15;
  reinterpret15_output_port_net <= b_16;
  clk_net <= clk_1;
  ce_net <= ce_1;
  mult0 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret0_output_port_net,
    b => reinterpret0_output_port_net_x0,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult0_p_net
  );
  mult1 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret1_output_port_net,
    b => reinterpret1_output_port_net_x0,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult1_p_net
  );
  mult2 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret2_output_port_net_x0,
    b => reinterpret2_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult2_p_net
  );
  mult3 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret3_output_port_net_x0,
    b => reinterpret3_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult3_p_net
  );
  mult4 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret4_output_port_net,
    b => reinterpret4_output_port_net_x0,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult4_p_net
  );
  mult5 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret5_output_port_net_x0,
    b => reinterpret5_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult5_p_net
  );
  mult6 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret6_output_port_net,
    b => reinterpret6_output_port_net_x0,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult6_p_net
  );
  mult7 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret7_output_port_net_x0,
    b => reinterpret7_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult7_p_net
  );
  mult8 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret8_output_port_net_x0,
    b => reinterpret8_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult8_p_net
  );
  mult9 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret9_output_port_net_x0,
    b => reinterpret9_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult9_p_net
  );
  mult10 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret10_output_port_net_x0,
    b => reinterpret10_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult10_p_net
  );
  mult11 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret11_output_port_net_x0,
    b => reinterpret11_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult11_p_net
  );
  mult12 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret12_output_port_net_x0,
    b => reinterpret12_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult12_p_net
  );
  mult13 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret13_output_port_net_x0,
    b => reinterpret13_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult13_p_net
  );
  mult14 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret14_output_port_net_x0,
    b => reinterpret14_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult14_p_net
  );
  mult15 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret15_output_port_net_x0,
    b => reinterpret15_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult15_p_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Vector Real Mult Im_2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_real_mult_im_2 is
  port (
    a_1 : in std_logic_vector( 16-1 downto 0 );
    b_1 : in std_logic_vector( 16-1 downto 0 );
    a_2 : in std_logic_vector( 16-1 downto 0 );
    a_3 : in std_logic_vector( 16-1 downto 0 );
    a_4 : in std_logic_vector( 16-1 downto 0 );
    a_5 : in std_logic_vector( 16-1 downto 0 );
    a_6 : in std_logic_vector( 16-1 downto 0 );
    a_7 : in std_logic_vector( 16-1 downto 0 );
    a_8 : in std_logic_vector( 16-1 downto 0 );
    a_9 : in std_logic_vector( 16-1 downto 0 );
    a_10 : in std_logic_vector( 16-1 downto 0 );
    a_11 : in std_logic_vector( 16-1 downto 0 );
    a_12 : in std_logic_vector( 16-1 downto 0 );
    a_13 : in std_logic_vector( 16-1 downto 0 );
    a_14 : in std_logic_vector( 16-1 downto 0 );
    a_15 : in std_logic_vector( 16-1 downto 0 );
    a_16 : in std_logic_vector( 16-1 downto 0 );
    b_2 : in std_logic_vector( 16-1 downto 0 );
    b_3 : in std_logic_vector( 16-1 downto 0 );
    b_4 : in std_logic_vector( 16-1 downto 0 );
    b_5 : in std_logic_vector( 16-1 downto 0 );
    b_6 : in std_logic_vector( 16-1 downto 0 );
    b_7 : in std_logic_vector( 16-1 downto 0 );
    b_8 : in std_logic_vector( 16-1 downto 0 );
    b_9 : in std_logic_vector( 16-1 downto 0 );
    b_10 : in std_logic_vector( 16-1 downto 0 );
    b_11 : in std_logic_vector( 16-1 downto 0 );
    b_12 : in std_logic_vector( 16-1 downto 0 );
    b_13 : in std_logic_vector( 16-1 downto 0 );
    b_14 : in std_logic_vector( 16-1 downto 0 );
    b_15 : in std_logic_vector( 16-1 downto 0 );
    b_16 : in std_logic_vector( 16-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    a_x_b_1 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_2 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_3 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_4 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_5 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_6 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_7 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_8 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_9 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_10 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_11 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_12 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_13 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_14 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_15 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_16 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_vector_real_mult_im_2;
architecture structural of psb3_0_vector_real_mult_im_2 is 
  signal reinterpret2_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal mult9_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal mult0_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult1_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal mult3_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mult6_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mult11_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult12_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal mult2_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal mult7_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult5_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult10_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult13_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult4_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult14_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult8_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult15_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal clk_net : std_logic;
  signal reinterpret14_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal ce_net : std_logic;
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
begin
  a_x_b_1 <= mult0_p_net;
  a_x_b_2 <= mult1_p_net;
  a_x_b_3 <= mult2_p_net;
  a_x_b_4 <= mult3_p_net;
  a_x_b_5 <= mult4_p_net;
  a_x_b_6 <= mult5_p_net;
  a_x_b_7 <= mult6_p_net;
  a_x_b_8 <= mult7_p_net;
  a_x_b_9 <= mult8_p_net;
  a_x_b_10 <= mult9_p_net;
  a_x_b_11 <= mult10_p_net;
  a_x_b_12 <= mult11_p_net;
  a_x_b_13 <= mult12_p_net;
  a_x_b_14 <= mult13_p_net;
  a_x_b_15 <= mult14_p_net;
  a_x_b_16 <= mult15_p_net;
  reinterpret0_output_port_net <= a_1;
  reinterpret0_output_port_net_x0 <= b_1;
  reinterpret1_output_port_net <= a_2;
  reinterpret2_output_port_net_x0 <= a_3;
  reinterpret3_output_port_net_x0 <= a_4;
  reinterpret4_output_port_net <= a_5;
  reinterpret5_output_port_net_x0 <= a_6;
  reinterpret6_output_port_net <= a_7;
  reinterpret7_output_port_net_x0 <= a_8;
  reinterpret8_output_port_net_x0 <= a_9;
  reinterpret9_output_port_net_x0 <= a_10;
  reinterpret10_output_port_net_x0 <= a_11;
  reinterpret11_output_port_net_x0 <= a_12;
  reinterpret12_output_port_net_x0 <= a_13;
  reinterpret13_output_port_net_x0 <= a_14;
  reinterpret14_output_port_net_x0 <= a_15;
  reinterpret15_output_port_net_x0 <= a_16;
  reinterpret1_output_port_net_x0 <= b_2;
  reinterpret2_output_port_net <= b_3;
  reinterpret3_output_port_net <= b_4;
  reinterpret4_output_port_net_x0 <= b_5;
  reinterpret5_output_port_net <= b_6;
  reinterpret6_output_port_net_x0 <= b_7;
  reinterpret7_output_port_net <= b_8;
  reinterpret8_output_port_net <= b_9;
  reinterpret9_output_port_net <= b_10;
  reinterpret10_output_port_net <= b_11;
  reinterpret11_output_port_net <= b_12;
  reinterpret12_output_port_net <= b_13;
  reinterpret13_output_port_net <= b_14;
  reinterpret14_output_port_net <= b_15;
  reinterpret15_output_port_net <= b_16;
  clk_net <= clk_1;
  ce_net <= ce_1;
  mult0 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret0_output_port_net,
    b => reinterpret0_output_port_net_x0,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult0_p_net
  );
  mult1 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret1_output_port_net,
    b => reinterpret1_output_port_net_x0,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult1_p_net
  );
  mult2 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret2_output_port_net_x0,
    b => reinterpret2_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult2_p_net
  );
  mult3 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret3_output_port_net_x0,
    b => reinterpret3_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult3_p_net
  );
  mult4 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret4_output_port_net,
    b => reinterpret4_output_port_net_x0,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult4_p_net
  );
  mult5 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret5_output_port_net_x0,
    b => reinterpret5_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult5_p_net
  );
  mult6 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret6_output_port_net,
    b => reinterpret6_output_port_net_x0,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult6_p_net
  );
  mult7 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret7_output_port_net_x0,
    b => reinterpret7_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult7_p_net
  );
  mult8 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret8_output_port_net_x0,
    b => reinterpret8_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult8_p_net
  );
  mult9 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret9_output_port_net_x0,
    b => reinterpret9_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult9_p_net
  );
  mult10 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret10_output_port_net_x0,
    b => reinterpret10_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult10_p_net
  );
  mult11 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret11_output_port_net_x0,
    b => reinterpret11_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult11_p_net
  );
  mult12 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret12_output_port_net_x0,
    b => reinterpret12_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult12_p_net
  );
  mult13 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret13_output_port_net_x0,
    b => reinterpret13_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult13_p_net
  );
  mult14 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret14_output_port_net_x0,
    b => reinterpret14_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult14_p_net
  );
  mult15 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret15_output_port_net_x0,
    b => reinterpret15_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult15_p_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Vector Real Mult Im_3
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_real_mult_im_3 is
  port (
    a_1 : in std_logic_vector( 16-1 downto 0 );
    b_1 : in std_logic_vector( 16-1 downto 0 );
    a_2 : in std_logic_vector( 16-1 downto 0 );
    a_3 : in std_logic_vector( 16-1 downto 0 );
    a_4 : in std_logic_vector( 16-1 downto 0 );
    a_5 : in std_logic_vector( 16-1 downto 0 );
    a_6 : in std_logic_vector( 16-1 downto 0 );
    a_7 : in std_logic_vector( 16-1 downto 0 );
    a_8 : in std_logic_vector( 16-1 downto 0 );
    a_9 : in std_logic_vector( 16-1 downto 0 );
    a_10 : in std_logic_vector( 16-1 downto 0 );
    a_11 : in std_logic_vector( 16-1 downto 0 );
    a_12 : in std_logic_vector( 16-1 downto 0 );
    a_13 : in std_logic_vector( 16-1 downto 0 );
    a_14 : in std_logic_vector( 16-1 downto 0 );
    a_15 : in std_logic_vector( 16-1 downto 0 );
    a_16 : in std_logic_vector( 16-1 downto 0 );
    b_2 : in std_logic_vector( 16-1 downto 0 );
    b_3 : in std_logic_vector( 16-1 downto 0 );
    b_4 : in std_logic_vector( 16-1 downto 0 );
    b_5 : in std_logic_vector( 16-1 downto 0 );
    b_6 : in std_logic_vector( 16-1 downto 0 );
    b_7 : in std_logic_vector( 16-1 downto 0 );
    b_8 : in std_logic_vector( 16-1 downto 0 );
    b_9 : in std_logic_vector( 16-1 downto 0 );
    b_10 : in std_logic_vector( 16-1 downto 0 );
    b_11 : in std_logic_vector( 16-1 downto 0 );
    b_12 : in std_logic_vector( 16-1 downto 0 );
    b_13 : in std_logic_vector( 16-1 downto 0 );
    b_14 : in std_logic_vector( 16-1 downto 0 );
    b_15 : in std_logic_vector( 16-1 downto 0 );
    b_16 : in std_logic_vector( 16-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    a_x_b_1 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_2 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_3 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_4 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_5 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_6 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_7 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_8 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_9 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_10 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_11 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_12 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_13 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_14 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_15 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_16 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_vector_real_mult_im_3;
architecture structural of psb3_0_vector_real_mult_im_3 is 
  signal mult13_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult8_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mult0_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult10_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mult1_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult6_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult5_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult3_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult9_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult12_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult2_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult4_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult11_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult7_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult14_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult15_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal clk_net : std_logic;
  signal reinterpret9_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal ce_net : std_logic;
  signal reinterpret1_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
begin
  a_x_b_1 <= mult0_p_net;
  a_x_b_2 <= mult1_p_net;
  a_x_b_3 <= mult2_p_net;
  a_x_b_4 <= mult3_p_net;
  a_x_b_5 <= mult4_p_net;
  a_x_b_6 <= mult5_p_net;
  a_x_b_7 <= mult6_p_net;
  a_x_b_8 <= mult7_p_net;
  a_x_b_9 <= mult8_p_net;
  a_x_b_10 <= mult9_p_net;
  a_x_b_11 <= mult10_p_net;
  a_x_b_12 <= mult11_p_net;
  a_x_b_13 <= mult12_p_net;
  a_x_b_14 <= mult13_p_net;
  a_x_b_15 <= mult14_p_net;
  a_x_b_16 <= mult15_p_net;
  reinterpret0_output_port_net <= a_1;
  reinterpret0_output_port_net_x0 <= b_1;
  reinterpret1_output_port_net <= a_2;
  reinterpret2_output_port_net_x0 <= a_3;
  reinterpret3_output_port_net_x0 <= a_4;
  reinterpret4_output_port_net <= a_5;
  reinterpret5_output_port_net_x0 <= a_6;
  reinterpret6_output_port_net <= a_7;
  reinterpret7_output_port_net_x0 <= a_8;
  reinterpret8_output_port_net_x0 <= a_9;
  reinterpret9_output_port_net_x0 <= a_10;
  reinterpret10_output_port_net_x0 <= a_11;
  reinterpret11_output_port_net_x0 <= a_12;
  reinterpret12_output_port_net_x0 <= a_13;
  reinterpret13_output_port_net_x0 <= a_14;
  reinterpret14_output_port_net_x0 <= a_15;
  reinterpret15_output_port_net_x0 <= a_16;
  reinterpret1_output_port_net_x0 <= b_2;
  reinterpret2_output_port_net <= b_3;
  reinterpret3_output_port_net <= b_4;
  reinterpret4_output_port_net_x0 <= b_5;
  reinterpret5_output_port_net <= b_6;
  reinterpret6_output_port_net_x0 <= b_7;
  reinterpret7_output_port_net <= b_8;
  reinterpret8_output_port_net <= b_9;
  reinterpret9_output_port_net <= b_10;
  reinterpret10_output_port_net <= b_11;
  reinterpret11_output_port_net <= b_12;
  reinterpret12_output_port_net <= b_13;
  reinterpret13_output_port_net <= b_14;
  reinterpret14_output_port_net <= b_15;
  reinterpret15_output_port_net <= b_16;
  clk_net <= clk_1;
  ce_net <= ce_1;
  mult0 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret0_output_port_net,
    b => reinterpret0_output_port_net_x0,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult0_p_net
  );
  mult1 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret1_output_port_net,
    b => reinterpret1_output_port_net_x0,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult1_p_net
  );
  mult2 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret2_output_port_net_x0,
    b => reinterpret2_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult2_p_net
  );
  mult3 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret3_output_port_net_x0,
    b => reinterpret3_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult3_p_net
  );
  mult4 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret4_output_port_net,
    b => reinterpret4_output_port_net_x0,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult4_p_net
  );
  mult5 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret5_output_port_net_x0,
    b => reinterpret5_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult5_p_net
  );
  mult6 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret6_output_port_net,
    b => reinterpret6_output_port_net_x0,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult6_p_net
  );
  mult7 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret7_output_port_net_x0,
    b => reinterpret7_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult7_p_net
  );
  mult8 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret8_output_port_net_x0,
    b => reinterpret8_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult8_p_net
  );
  mult9 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret9_output_port_net_x0,
    b => reinterpret9_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult9_p_net
  );
  mult10 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret10_output_port_net_x0,
    b => reinterpret10_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult10_p_net
  );
  mult11 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret11_output_port_net_x0,
    b => reinterpret11_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult11_p_net
  );
  mult12 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret12_output_port_net_x0,
    b => reinterpret12_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult12_p_net
  );
  mult13 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret13_output_port_net_x0,
    b => reinterpret13_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult13_p_net
  );
  mult14 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret14_output_port_net_x0,
    b => reinterpret14_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult14_p_net
  );
  mult15 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret15_output_port_net_x0,
    b => reinterpret15_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult15_p_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Vector Real Mult Im_4
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_real_mult_im_4 is
  port (
    a_1 : in std_logic_vector( 16-1 downto 0 );
    b_1 : in std_logic_vector( 16-1 downto 0 );
    a_2 : in std_logic_vector( 16-1 downto 0 );
    a_3 : in std_logic_vector( 16-1 downto 0 );
    a_4 : in std_logic_vector( 16-1 downto 0 );
    a_5 : in std_logic_vector( 16-1 downto 0 );
    a_6 : in std_logic_vector( 16-1 downto 0 );
    a_7 : in std_logic_vector( 16-1 downto 0 );
    a_8 : in std_logic_vector( 16-1 downto 0 );
    a_9 : in std_logic_vector( 16-1 downto 0 );
    a_10 : in std_logic_vector( 16-1 downto 0 );
    a_11 : in std_logic_vector( 16-1 downto 0 );
    a_12 : in std_logic_vector( 16-1 downto 0 );
    a_13 : in std_logic_vector( 16-1 downto 0 );
    a_14 : in std_logic_vector( 16-1 downto 0 );
    a_15 : in std_logic_vector( 16-1 downto 0 );
    a_16 : in std_logic_vector( 16-1 downto 0 );
    b_2 : in std_logic_vector( 16-1 downto 0 );
    b_3 : in std_logic_vector( 16-1 downto 0 );
    b_4 : in std_logic_vector( 16-1 downto 0 );
    b_5 : in std_logic_vector( 16-1 downto 0 );
    b_6 : in std_logic_vector( 16-1 downto 0 );
    b_7 : in std_logic_vector( 16-1 downto 0 );
    b_8 : in std_logic_vector( 16-1 downto 0 );
    b_9 : in std_logic_vector( 16-1 downto 0 );
    b_10 : in std_logic_vector( 16-1 downto 0 );
    b_11 : in std_logic_vector( 16-1 downto 0 );
    b_12 : in std_logic_vector( 16-1 downto 0 );
    b_13 : in std_logic_vector( 16-1 downto 0 );
    b_14 : in std_logic_vector( 16-1 downto 0 );
    b_15 : in std_logic_vector( 16-1 downto 0 );
    b_16 : in std_logic_vector( 16-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    a_x_b_1 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_2 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_3 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_4 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_5 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_6 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_7 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_8 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_9 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_10 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_11 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_12 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_13 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_14 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_15 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_16 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_vector_real_mult_im_4;
architecture structural of psb3_0_vector_real_mult_im_4 is 
  signal mult4_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult2_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult3_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult5_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult6_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult7_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult1_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult8_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult0_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal mult10_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal mult15_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal mult12_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal mult11_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal mult9_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal mult13_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult14_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal ce_net : std_logic;
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal clk_net : std_logic;
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
begin
  a_x_b_1 <= mult0_p_net;
  a_x_b_2 <= mult1_p_net;
  a_x_b_3 <= mult2_p_net;
  a_x_b_4 <= mult3_p_net;
  a_x_b_5 <= mult4_p_net;
  a_x_b_6 <= mult5_p_net;
  a_x_b_7 <= mult6_p_net;
  a_x_b_8 <= mult7_p_net;
  a_x_b_9 <= mult8_p_net;
  a_x_b_10 <= mult9_p_net;
  a_x_b_11 <= mult10_p_net;
  a_x_b_12 <= mult11_p_net;
  a_x_b_13 <= mult12_p_net;
  a_x_b_14 <= mult13_p_net;
  a_x_b_15 <= mult14_p_net;
  a_x_b_16 <= mult15_p_net;
  reinterpret0_output_port_net <= a_1;
  reinterpret0_output_port_net_x0 <= b_1;
  reinterpret1_output_port_net <= a_2;
  reinterpret2_output_port_net_x0 <= a_3;
  reinterpret3_output_port_net_x0 <= a_4;
  reinterpret4_output_port_net <= a_5;
  reinterpret5_output_port_net_x0 <= a_6;
  reinterpret6_output_port_net <= a_7;
  reinterpret7_output_port_net_x0 <= a_8;
  reinterpret8_output_port_net_x0 <= a_9;
  reinterpret9_output_port_net_x0 <= a_10;
  reinterpret10_output_port_net_x0 <= a_11;
  reinterpret11_output_port_net_x0 <= a_12;
  reinterpret12_output_port_net_x0 <= a_13;
  reinterpret13_output_port_net_x0 <= a_14;
  reinterpret14_output_port_net_x0 <= a_15;
  reinterpret15_output_port_net_x0 <= a_16;
  reinterpret1_output_port_net_x0 <= b_2;
  reinterpret2_output_port_net <= b_3;
  reinterpret3_output_port_net <= b_4;
  reinterpret4_output_port_net_x0 <= b_5;
  reinterpret5_output_port_net <= b_6;
  reinterpret6_output_port_net_x0 <= b_7;
  reinterpret7_output_port_net <= b_8;
  reinterpret8_output_port_net <= b_9;
  reinterpret9_output_port_net <= b_10;
  reinterpret10_output_port_net <= b_11;
  reinterpret11_output_port_net <= b_12;
  reinterpret12_output_port_net <= b_13;
  reinterpret13_output_port_net <= b_14;
  reinterpret14_output_port_net <= b_15;
  reinterpret15_output_port_net <= b_16;
  clk_net <= clk_1;
  ce_net <= ce_1;
  mult0 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret0_output_port_net,
    b => reinterpret0_output_port_net_x0,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult0_p_net
  );
  mult1 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret1_output_port_net,
    b => reinterpret1_output_port_net_x0,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult1_p_net
  );
  mult2 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret2_output_port_net_x0,
    b => reinterpret2_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult2_p_net
  );
  mult3 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret3_output_port_net_x0,
    b => reinterpret3_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult3_p_net
  );
  mult4 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret4_output_port_net,
    b => reinterpret4_output_port_net_x0,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult4_p_net
  );
  mult5 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret5_output_port_net_x0,
    b => reinterpret5_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult5_p_net
  );
  mult6 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret6_output_port_net,
    b => reinterpret6_output_port_net_x0,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult6_p_net
  );
  mult7 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret7_output_port_net_x0,
    b => reinterpret7_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult7_p_net
  );
  mult8 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret8_output_port_net_x0,
    b => reinterpret8_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult8_p_net
  );
  mult9 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret9_output_port_net_x0,
    b => reinterpret9_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult9_p_net
  );
  mult10 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret10_output_port_net_x0,
    b => reinterpret10_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult10_p_net
  );
  mult11 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret11_output_port_net_x0,
    b => reinterpret11_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult11_p_net
  );
  mult12 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret12_output_port_net_x0,
    b => reinterpret12_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult12_p_net
  );
  mult13 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret13_output_port_net_x0,
    b => reinterpret13_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult13_p_net
  );
  mult14 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret14_output_port_net_x0,
    b => reinterpret14_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult14_p_net
  );
  mult15 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret15_output_port_net_x0,
    b => reinterpret15_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult15_p_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Vector Real Mult Re_1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_real_mult_re_1 is
  port (
    a_1 : in std_logic_vector( 16-1 downto 0 );
    b_1 : in std_logic_vector( 16-1 downto 0 );
    a_2 : in std_logic_vector( 16-1 downto 0 );
    a_3 : in std_logic_vector( 16-1 downto 0 );
    a_4 : in std_logic_vector( 16-1 downto 0 );
    a_5 : in std_logic_vector( 16-1 downto 0 );
    a_6 : in std_logic_vector( 16-1 downto 0 );
    a_7 : in std_logic_vector( 16-1 downto 0 );
    a_8 : in std_logic_vector( 16-1 downto 0 );
    a_9 : in std_logic_vector( 16-1 downto 0 );
    a_10 : in std_logic_vector( 16-1 downto 0 );
    a_11 : in std_logic_vector( 16-1 downto 0 );
    a_12 : in std_logic_vector( 16-1 downto 0 );
    a_13 : in std_logic_vector( 16-1 downto 0 );
    a_14 : in std_logic_vector( 16-1 downto 0 );
    a_15 : in std_logic_vector( 16-1 downto 0 );
    a_16 : in std_logic_vector( 16-1 downto 0 );
    b_2 : in std_logic_vector( 16-1 downto 0 );
    b_3 : in std_logic_vector( 16-1 downto 0 );
    b_4 : in std_logic_vector( 16-1 downto 0 );
    b_5 : in std_logic_vector( 16-1 downto 0 );
    b_6 : in std_logic_vector( 16-1 downto 0 );
    b_7 : in std_logic_vector( 16-1 downto 0 );
    b_8 : in std_logic_vector( 16-1 downto 0 );
    b_9 : in std_logic_vector( 16-1 downto 0 );
    b_10 : in std_logic_vector( 16-1 downto 0 );
    b_11 : in std_logic_vector( 16-1 downto 0 );
    b_12 : in std_logic_vector( 16-1 downto 0 );
    b_13 : in std_logic_vector( 16-1 downto 0 );
    b_14 : in std_logic_vector( 16-1 downto 0 );
    b_15 : in std_logic_vector( 16-1 downto 0 );
    b_16 : in std_logic_vector( 16-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    a_x_b_1 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_2 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_3 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_4 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_5 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_6 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_7 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_8 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_9 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_10 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_11 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_12 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_13 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_14 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_15 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_16 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_vector_real_mult_re_1;
architecture structural of psb3_0_vector_real_mult_re_1 is 
  signal reinterpret8_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal mult3_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal mult6_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult12_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult7_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult13_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal mult14_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal mult4_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult9_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult11_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult15_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mult1_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult2_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal mult5_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal mult0_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult8_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult10_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal ce_net : std_logic;
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal clk_net : std_logic;
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
begin
  a_x_b_1 <= mult0_p_net;
  a_x_b_2 <= mult1_p_net;
  a_x_b_3 <= mult2_p_net;
  a_x_b_4 <= mult3_p_net;
  a_x_b_5 <= mult4_p_net;
  a_x_b_6 <= mult5_p_net;
  a_x_b_7 <= mult6_p_net;
  a_x_b_8 <= mult7_p_net;
  a_x_b_9 <= mult8_p_net;
  a_x_b_10 <= mult9_p_net;
  a_x_b_11 <= mult10_p_net;
  a_x_b_12 <= mult11_p_net;
  a_x_b_13 <= mult12_p_net;
  a_x_b_14 <= mult13_p_net;
  a_x_b_15 <= mult14_p_net;
  a_x_b_16 <= mult15_p_net;
  reinterpret0_output_port_net <= a_1;
  reinterpret0_output_port_net_x0 <= b_1;
  reinterpret1_output_port_net <= a_2;
  reinterpret2_output_port_net_x0 <= a_3;
  reinterpret3_output_port_net_x0 <= a_4;
  reinterpret4_output_port_net <= a_5;
  reinterpret5_output_port_net_x0 <= a_6;
  reinterpret6_output_port_net <= a_7;
  reinterpret7_output_port_net_x0 <= a_8;
  reinterpret8_output_port_net_x0 <= a_9;
  reinterpret9_output_port_net_x0 <= a_10;
  reinterpret10_output_port_net_x0 <= a_11;
  reinterpret11_output_port_net_x0 <= a_12;
  reinterpret12_output_port_net_x0 <= a_13;
  reinterpret13_output_port_net_x0 <= a_14;
  reinterpret14_output_port_net_x0 <= a_15;
  reinterpret15_output_port_net_x0 <= a_16;
  reinterpret1_output_port_net_x0 <= b_2;
  reinterpret2_output_port_net <= b_3;
  reinterpret3_output_port_net <= b_4;
  reinterpret4_output_port_net_x0 <= b_5;
  reinterpret5_output_port_net <= b_6;
  reinterpret6_output_port_net_x0 <= b_7;
  reinterpret7_output_port_net <= b_8;
  reinterpret8_output_port_net <= b_9;
  reinterpret9_output_port_net <= b_10;
  reinterpret10_output_port_net <= b_11;
  reinterpret11_output_port_net <= b_12;
  reinterpret12_output_port_net <= b_13;
  reinterpret13_output_port_net <= b_14;
  reinterpret14_output_port_net <= b_15;
  reinterpret15_output_port_net <= b_16;
  clk_net <= clk_1;
  ce_net <= ce_1;
  mult0 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret0_output_port_net,
    b => reinterpret0_output_port_net_x0,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult0_p_net
  );
  mult1 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret1_output_port_net,
    b => reinterpret1_output_port_net_x0,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult1_p_net
  );
  mult2 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret2_output_port_net_x0,
    b => reinterpret2_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult2_p_net
  );
  mult3 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret3_output_port_net_x0,
    b => reinterpret3_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult3_p_net
  );
  mult4 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret4_output_port_net,
    b => reinterpret4_output_port_net_x0,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult4_p_net
  );
  mult5 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret5_output_port_net_x0,
    b => reinterpret5_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult5_p_net
  );
  mult6 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret6_output_port_net,
    b => reinterpret6_output_port_net_x0,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult6_p_net
  );
  mult7 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret7_output_port_net_x0,
    b => reinterpret7_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult7_p_net
  );
  mult8 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret8_output_port_net_x0,
    b => reinterpret8_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult8_p_net
  );
  mult9 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret9_output_port_net_x0,
    b => reinterpret9_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult9_p_net
  );
  mult10 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret10_output_port_net_x0,
    b => reinterpret10_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult10_p_net
  );
  mult11 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret11_output_port_net_x0,
    b => reinterpret11_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult11_p_net
  );
  mult12 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret12_output_port_net_x0,
    b => reinterpret12_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult12_p_net
  );
  mult13 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret13_output_port_net_x0,
    b => reinterpret13_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult13_p_net
  );
  mult14 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret14_output_port_net_x0,
    b => reinterpret14_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult14_p_net
  );
  mult15 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret15_output_port_net_x0,
    b => reinterpret15_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult15_p_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Vector Real Mult Re_2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_real_mult_re_2 is
  port (
    a_1 : in std_logic_vector( 16-1 downto 0 );
    b_1 : in std_logic_vector( 16-1 downto 0 );
    a_2 : in std_logic_vector( 16-1 downto 0 );
    a_3 : in std_logic_vector( 16-1 downto 0 );
    a_4 : in std_logic_vector( 16-1 downto 0 );
    a_5 : in std_logic_vector( 16-1 downto 0 );
    a_6 : in std_logic_vector( 16-1 downto 0 );
    a_7 : in std_logic_vector( 16-1 downto 0 );
    a_8 : in std_logic_vector( 16-1 downto 0 );
    a_9 : in std_logic_vector( 16-1 downto 0 );
    a_10 : in std_logic_vector( 16-1 downto 0 );
    a_11 : in std_logic_vector( 16-1 downto 0 );
    a_12 : in std_logic_vector( 16-1 downto 0 );
    a_13 : in std_logic_vector( 16-1 downto 0 );
    a_14 : in std_logic_vector( 16-1 downto 0 );
    a_15 : in std_logic_vector( 16-1 downto 0 );
    a_16 : in std_logic_vector( 16-1 downto 0 );
    b_2 : in std_logic_vector( 16-1 downto 0 );
    b_3 : in std_logic_vector( 16-1 downto 0 );
    b_4 : in std_logic_vector( 16-1 downto 0 );
    b_5 : in std_logic_vector( 16-1 downto 0 );
    b_6 : in std_logic_vector( 16-1 downto 0 );
    b_7 : in std_logic_vector( 16-1 downto 0 );
    b_8 : in std_logic_vector( 16-1 downto 0 );
    b_9 : in std_logic_vector( 16-1 downto 0 );
    b_10 : in std_logic_vector( 16-1 downto 0 );
    b_11 : in std_logic_vector( 16-1 downto 0 );
    b_12 : in std_logic_vector( 16-1 downto 0 );
    b_13 : in std_logic_vector( 16-1 downto 0 );
    b_14 : in std_logic_vector( 16-1 downto 0 );
    b_15 : in std_logic_vector( 16-1 downto 0 );
    b_16 : in std_logic_vector( 16-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    a_x_b_1 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_2 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_3 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_4 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_5 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_6 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_7 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_8 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_9 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_10 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_11 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_12 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_13 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_14 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_15 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_16 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_vector_real_mult_re_2;
architecture structural of psb3_0_vector_real_mult_re_2 is 
  signal mult13_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult5_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult15_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal mult10_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal mult2_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult9_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult8_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult12_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult6_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult14_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult1_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult4_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult7_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult0_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult3_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult11_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal ce_net : std_logic;
  signal reinterpret11_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal clk_net : std_logic;
  signal reinterpret3_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
begin
  a_x_b_1 <= mult0_p_net;
  a_x_b_2 <= mult1_p_net;
  a_x_b_3 <= mult2_p_net;
  a_x_b_4 <= mult3_p_net;
  a_x_b_5 <= mult4_p_net;
  a_x_b_6 <= mult5_p_net;
  a_x_b_7 <= mult6_p_net;
  a_x_b_8 <= mult7_p_net;
  a_x_b_9 <= mult8_p_net;
  a_x_b_10 <= mult9_p_net;
  a_x_b_11 <= mult10_p_net;
  a_x_b_12 <= mult11_p_net;
  a_x_b_13 <= mult12_p_net;
  a_x_b_14 <= mult13_p_net;
  a_x_b_15 <= mult14_p_net;
  a_x_b_16 <= mult15_p_net;
  reinterpret0_output_port_net <= a_1;
  reinterpret0_output_port_net_x0 <= b_1;
  reinterpret1_output_port_net <= a_2;
  reinterpret2_output_port_net_x0 <= a_3;
  reinterpret3_output_port_net_x0 <= a_4;
  reinterpret4_output_port_net <= a_5;
  reinterpret5_output_port_net_x0 <= a_6;
  reinterpret6_output_port_net <= a_7;
  reinterpret7_output_port_net_x0 <= a_8;
  reinterpret8_output_port_net_x0 <= a_9;
  reinterpret9_output_port_net_x0 <= a_10;
  reinterpret10_output_port_net_x0 <= a_11;
  reinterpret11_output_port_net_x0 <= a_12;
  reinterpret12_output_port_net_x0 <= a_13;
  reinterpret13_output_port_net_x0 <= a_14;
  reinterpret14_output_port_net_x0 <= a_15;
  reinterpret15_output_port_net_x0 <= a_16;
  reinterpret1_output_port_net_x0 <= b_2;
  reinterpret2_output_port_net <= b_3;
  reinterpret3_output_port_net <= b_4;
  reinterpret4_output_port_net_x0 <= b_5;
  reinterpret5_output_port_net <= b_6;
  reinterpret6_output_port_net_x0 <= b_7;
  reinterpret7_output_port_net <= b_8;
  reinterpret8_output_port_net <= b_9;
  reinterpret9_output_port_net <= b_10;
  reinterpret10_output_port_net <= b_11;
  reinterpret11_output_port_net <= b_12;
  reinterpret12_output_port_net <= b_13;
  reinterpret13_output_port_net <= b_14;
  reinterpret14_output_port_net <= b_15;
  reinterpret15_output_port_net <= b_16;
  clk_net <= clk_1;
  ce_net <= ce_1;
  mult0 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret0_output_port_net,
    b => reinterpret0_output_port_net_x0,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult0_p_net
  );
  mult1 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret1_output_port_net,
    b => reinterpret1_output_port_net_x0,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult1_p_net
  );
  mult2 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret2_output_port_net_x0,
    b => reinterpret2_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult2_p_net
  );
  mult3 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret3_output_port_net_x0,
    b => reinterpret3_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult3_p_net
  );
  mult4 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret4_output_port_net,
    b => reinterpret4_output_port_net_x0,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult4_p_net
  );
  mult5 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret5_output_port_net_x0,
    b => reinterpret5_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult5_p_net
  );
  mult6 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret6_output_port_net,
    b => reinterpret6_output_port_net_x0,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult6_p_net
  );
  mult7 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret7_output_port_net_x0,
    b => reinterpret7_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult7_p_net
  );
  mult8 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret8_output_port_net_x0,
    b => reinterpret8_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult8_p_net
  );
  mult9 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret9_output_port_net_x0,
    b => reinterpret9_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult9_p_net
  );
  mult10 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret10_output_port_net_x0,
    b => reinterpret10_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult10_p_net
  );
  mult11 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret11_output_port_net_x0,
    b => reinterpret11_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult11_p_net
  );
  mult12 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret12_output_port_net_x0,
    b => reinterpret12_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult12_p_net
  );
  mult13 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret13_output_port_net_x0,
    b => reinterpret13_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult13_p_net
  );
  mult14 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret14_output_port_net_x0,
    b => reinterpret14_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult14_p_net
  );
  mult15 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret15_output_port_net_x0,
    b => reinterpret15_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult15_p_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Vector Real Mult Re_3
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_real_mult_re_3 is
  port (
    a_1 : in std_logic_vector( 16-1 downto 0 );
    b_1 : in std_logic_vector( 16-1 downto 0 );
    a_2 : in std_logic_vector( 16-1 downto 0 );
    a_3 : in std_logic_vector( 16-1 downto 0 );
    a_4 : in std_logic_vector( 16-1 downto 0 );
    a_5 : in std_logic_vector( 16-1 downto 0 );
    a_6 : in std_logic_vector( 16-1 downto 0 );
    a_7 : in std_logic_vector( 16-1 downto 0 );
    a_8 : in std_logic_vector( 16-1 downto 0 );
    a_9 : in std_logic_vector( 16-1 downto 0 );
    a_10 : in std_logic_vector( 16-1 downto 0 );
    a_11 : in std_logic_vector( 16-1 downto 0 );
    a_12 : in std_logic_vector( 16-1 downto 0 );
    a_13 : in std_logic_vector( 16-1 downto 0 );
    a_14 : in std_logic_vector( 16-1 downto 0 );
    a_15 : in std_logic_vector( 16-1 downto 0 );
    a_16 : in std_logic_vector( 16-1 downto 0 );
    b_2 : in std_logic_vector( 16-1 downto 0 );
    b_3 : in std_logic_vector( 16-1 downto 0 );
    b_4 : in std_logic_vector( 16-1 downto 0 );
    b_5 : in std_logic_vector( 16-1 downto 0 );
    b_6 : in std_logic_vector( 16-1 downto 0 );
    b_7 : in std_logic_vector( 16-1 downto 0 );
    b_8 : in std_logic_vector( 16-1 downto 0 );
    b_9 : in std_logic_vector( 16-1 downto 0 );
    b_10 : in std_logic_vector( 16-1 downto 0 );
    b_11 : in std_logic_vector( 16-1 downto 0 );
    b_12 : in std_logic_vector( 16-1 downto 0 );
    b_13 : in std_logic_vector( 16-1 downto 0 );
    b_14 : in std_logic_vector( 16-1 downto 0 );
    b_15 : in std_logic_vector( 16-1 downto 0 );
    b_16 : in std_logic_vector( 16-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    a_x_b_1 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_2 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_3 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_4 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_5 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_6 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_7 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_8 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_9 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_10 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_11 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_12 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_13 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_14 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_15 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_16 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_vector_real_mult_re_3;
architecture structural of psb3_0_vector_real_mult_re_3 is 
  signal reinterpret9_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal mult14_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mult11_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal mult8_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult9_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal mult12_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult10_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult15_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult13_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal mult5_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult7_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult6_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult0_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult1_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult2_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult3_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult4_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal ce_net : std_logic;
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal clk_net : std_logic;
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
begin
  a_x_b_1 <= mult0_p_net;
  a_x_b_2 <= mult1_p_net;
  a_x_b_3 <= mult2_p_net;
  a_x_b_4 <= mult3_p_net;
  a_x_b_5 <= mult4_p_net;
  a_x_b_6 <= mult5_p_net;
  a_x_b_7 <= mult6_p_net;
  a_x_b_8 <= mult7_p_net;
  a_x_b_9 <= mult8_p_net;
  a_x_b_10 <= mult9_p_net;
  a_x_b_11 <= mult10_p_net;
  a_x_b_12 <= mult11_p_net;
  a_x_b_13 <= mult12_p_net;
  a_x_b_14 <= mult13_p_net;
  a_x_b_15 <= mult14_p_net;
  a_x_b_16 <= mult15_p_net;
  reinterpret0_output_port_net <= a_1;
  reinterpret0_output_port_net_x0 <= b_1;
  reinterpret1_output_port_net <= a_2;
  reinterpret2_output_port_net_x0 <= a_3;
  reinterpret3_output_port_net_x0 <= a_4;
  reinterpret4_output_port_net <= a_5;
  reinterpret5_output_port_net_x0 <= a_6;
  reinterpret6_output_port_net <= a_7;
  reinterpret7_output_port_net_x0 <= a_8;
  reinterpret8_output_port_net_x0 <= a_9;
  reinterpret9_output_port_net_x0 <= a_10;
  reinterpret10_output_port_net_x0 <= a_11;
  reinterpret11_output_port_net_x0 <= a_12;
  reinterpret12_output_port_net_x0 <= a_13;
  reinterpret13_output_port_net_x0 <= a_14;
  reinterpret14_output_port_net_x0 <= a_15;
  reinterpret15_output_port_net_x0 <= a_16;
  reinterpret1_output_port_net_x0 <= b_2;
  reinterpret2_output_port_net <= b_3;
  reinterpret3_output_port_net <= b_4;
  reinterpret4_output_port_net_x0 <= b_5;
  reinterpret5_output_port_net <= b_6;
  reinterpret6_output_port_net_x0 <= b_7;
  reinterpret7_output_port_net <= b_8;
  reinterpret8_output_port_net <= b_9;
  reinterpret9_output_port_net <= b_10;
  reinterpret10_output_port_net <= b_11;
  reinterpret11_output_port_net <= b_12;
  reinterpret12_output_port_net <= b_13;
  reinterpret13_output_port_net <= b_14;
  reinterpret14_output_port_net <= b_15;
  reinterpret15_output_port_net <= b_16;
  clk_net <= clk_1;
  ce_net <= ce_1;
  mult0 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret0_output_port_net,
    b => reinterpret0_output_port_net_x0,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult0_p_net
  );
  mult1 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret1_output_port_net,
    b => reinterpret1_output_port_net_x0,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult1_p_net
  );
  mult2 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret2_output_port_net_x0,
    b => reinterpret2_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult2_p_net
  );
  mult3 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret3_output_port_net_x0,
    b => reinterpret3_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult3_p_net
  );
  mult4 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret4_output_port_net,
    b => reinterpret4_output_port_net_x0,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult4_p_net
  );
  mult5 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret5_output_port_net_x0,
    b => reinterpret5_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult5_p_net
  );
  mult6 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret6_output_port_net,
    b => reinterpret6_output_port_net_x0,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult6_p_net
  );
  mult7 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret7_output_port_net_x0,
    b => reinterpret7_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult7_p_net
  );
  mult8 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret8_output_port_net_x0,
    b => reinterpret8_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult8_p_net
  );
  mult9 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret9_output_port_net_x0,
    b => reinterpret9_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult9_p_net
  );
  mult10 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret10_output_port_net_x0,
    b => reinterpret10_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult10_p_net
  );
  mult11 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret11_output_port_net_x0,
    b => reinterpret11_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult11_p_net
  );
  mult12 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret12_output_port_net_x0,
    b => reinterpret12_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult12_p_net
  );
  mult13 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret13_output_port_net_x0,
    b => reinterpret13_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult13_p_net
  );
  mult14 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret14_output_port_net_x0,
    b => reinterpret14_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult14_p_net
  );
  mult15 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret15_output_port_net_x0,
    b => reinterpret15_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult15_p_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Vector Real Mult Re_4
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_real_mult_re_4 is
  port (
    a_1 : in std_logic_vector( 16-1 downto 0 );
    b_1 : in std_logic_vector( 16-1 downto 0 );
    a_2 : in std_logic_vector( 16-1 downto 0 );
    a_3 : in std_logic_vector( 16-1 downto 0 );
    a_4 : in std_logic_vector( 16-1 downto 0 );
    a_5 : in std_logic_vector( 16-1 downto 0 );
    a_6 : in std_logic_vector( 16-1 downto 0 );
    a_7 : in std_logic_vector( 16-1 downto 0 );
    a_8 : in std_logic_vector( 16-1 downto 0 );
    a_9 : in std_logic_vector( 16-1 downto 0 );
    a_10 : in std_logic_vector( 16-1 downto 0 );
    a_11 : in std_logic_vector( 16-1 downto 0 );
    a_12 : in std_logic_vector( 16-1 downto 0 );
    a_13 : in std_logic_vector( 16-1 downto 0 );
    a_14 : in std_logic_vector( 16-1 downto 0 );
    a_15 : in std_logic_vector( 16-1 downto 0 );
    a_16 : in std_logic_vector( 16-1 downto 0 );
    b_2 : in std_logic_vector( 16-1 downto 0 );
    b_3 : in std_logic_vector( 16-1 downto 0 );
    b_4 : in std_logic_vector( 16-1 downto 0 );
    b_5 : in std_logic_vector( 16-1 downto 0 );
    b_6 : in std_logic_vector( 16-1 downto 0 );
    b_7 : in std_logic_vector( 16-1 downto 0 );
    b_8 : in std_logic_vector( 16-1 downto 0 );
    b_9 : in std_logic_vector( 16-1 downto 0 );
    b_10 : in std_logic_vector( 16-1 downto 0 );
    b_11 : in std_logic_vector( 16-1 downto 0 );
    b_12 : in std_logic_vector( 16-1 downto 0 );
    b_13 : in std_logic_vector( 16-1 downto 0 );
    b_14 : in std_logic_vector( 16-1 downto 0 );
    b_15 : in std_logic_vector( 16-1 downto 0 );
    b_16 : in std_logic_vector( 16-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    a_x_b_1 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_2 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_3 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_4 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_5 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_6 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_7 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_8 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_9 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_10 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_11 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_12 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_13 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_14 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_15 : out std_logic_vector( 16-1 downto 0 );
    a_x_b_16 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_vector_real_mult_re_4;
architecture structural of psb3_0_vector_real_mult_re_4 is 
  signal mult1_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mult6_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mult13_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal mult4_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult14_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal mult5_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult15_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult10_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal mult3_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult0_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mult7_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal mult12_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult2_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult8_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult9_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal mult11_p_net : std_logic_vector( 16-1 downto 0 );
  signal clk_net : std_logic;
  signal ce_net : std_logic;
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
begin
  a_x_b_1 <= mult0_p_net;
  a_x_b_2 <= mult1_p_net;
  a_x_b_3 <= mult2_p_net;
  a_x_b_4 <= mult3_p_net;
  a_x_b_5 <= mult4_p_net;
  a_x_b_6 <= mult5_p_net;
  a_x_b_7 <= mult6_p_net;
  a_x_b_8 <= mult7_p_net;
  a_x_b_9 <= mult8_p_net;
  a_x_b_10 <= mult9_p_net;
  a_x_b_11 <= mult10_p_net;
  a_x_b_12 <= mult11_p_net;
  a_x_b_13 <= mult12_p_net;
  a_x_b_14 <= mult13_p_net;
  a_x_b_15 <= mult14_p_net;
  a_x_b_16 <= mult15_p_net;
  reinterpret0_output_port_net <= a_1;
  reinterpret0_output_port_net_x0 <= b_1;
  reinterpret1_output_port_net <= a_2;
  reinterpret2_output_port_net_x0 <= a_3;
  reinterpret3_output_port_net_x0 <= a_4;
  reinterpret4_output_port_net <= a_5;
  reinterpret5_output_port_net_x0 <= a_6;
  reinterpret6_output_port_net <= a_7;
  reinterpret7_output_port_net_x0 <= a_8;
  reinterpret8_output_port_net_x0 <= a_9;
  reinterpret9_output_port_net_x0 <= a_10;
  reinterpret10_output_port_net_x0 <= a_11;
  reinterpret11_output_port_net_x0 <= a_12;
  reinterpret12_output_port_net_x0 <= a_13;
  reinterpret13_output_port_net_x0 <= a_14;
  reinterpret14_output_port_net_x0 <= a_15;
  reinterpret15_output_port_net_x0 <= a_16;
  reinterpret1_output_port_net_x0 <= b_2;
  reinterpret2_output_port_net <= b_3;
  reinterpret3_output_port_net <= b_4;
  reinterpret4_output_port_net_x0 <= b_5;
  reinterpret5_output_port_net <= b_6;
  reinterpret6_output_port_net_x0 <= b_7;
  reinterpret7_output_port_net <= b_8;
  reinterpret8_output_port_net <= b_9;
  reinterpret9_output_port_net <= b_10;
  reinterpret10_output_port_net <= b_11;
  reinterpret11_output_port_net <= b_12;
  reinterpret12_output_port_net <= b_13;
  reinterpret13_output_port_net <= b_14;
  reinterpret14_output_port_net <= b_15;
  reinterpret15_output_port_net <= b_16;
  clk_net <= clk_1;
  ce_net <= ce_1;
  mult0 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret0_output_port_net,
    b => reinterpret0_output_port_net_x0,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult0_p_net
  );
  mult1 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret1_output_port_net,
    b => reinterpret1_output_port_net_x0,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult1_p_net
  );
  mult2 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret2_output_port_net_x0,
    b => reinterpret2_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult2_p_net
  );
  mult3 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret3_output_port_net_x0,
    b => reinterpret3_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult3_p_net
  );
  mult4 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret4_output_port_net,
    b => reinterpret4_output_port_net_x0,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult4_p_net
  );
  mult5 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret5_output_port_net_x0,
    b => reinterpret5_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult5_p_net
  );
  mult6 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret6_output_port_net,
    b => reinterpret6_output_port_net_x0,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult6_p_net
  );
  mult7 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret7_output_port_net_x0,
    b => reinterpret7_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult7_p_net
  );
  mult8 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret8_output_port_net_x0,
    b => reinterpret8_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult8_p_net
  );
  mult9 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret9_output_port_net_x0,
    b => reinterpret9_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult9_p_net
  );
  mult10 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret10_output_port_net_x0,
    b => reinterpret10_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult10_p_net
  );
  mult11 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret11_output_port_net_x0,
    b => reinterpret11_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult11_p_net
  );
  mult12 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret12_output_port_net_x0,
    b => reinterpret12_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult12_p_net
  );
  mult13 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret13_output_port_net_x0,
    b => reinterpret13_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult13_p_net
  );
  mult14 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret14_output_port_net_x0,
    b => reinterpret14_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult14_p_net
  );
  mult15 : entity xil_defaultlib.psb3_0_xlmult 
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 15,
    a_width => 16,
    b_arith => xlSigned,
    b_bin_pt => 15,
    b_width => 16,
    c_a_type => 0,
    c_a_width => 16,
    c_b_type => 0,
    c_b_width => 16,
    c_baat => 16,
    c_output_width => 32,
    c_type => 0,
    core_name0 => "psb3_0_mult_gen_v12_0_i0",
    extra_registers => 2,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 15,
    p_width => 16,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => reinterpret15_output_port_net_x0,
    b => reinterpret15_output_port_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult15_p_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Vector Reinterpret1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_reinterpret1 is
  port (
    in_1 : in std_logic_vector( 16-1 downto 0 );
    in_2 : in std_logic_vector( 16-1 downto 0 );
    in_3 : in std_logic_vector( 16-1 downto 0 );
    in_4 : in std_logic_vector( 16-1 downto 0 );
    in_5 : in std_logic_vector( 16-1 downto 0 );
    in_6 : in std_logic_vector( 16-1 downto 0 );
    in_7 : in std_logic_vector( 16-1 downto 0 );
    in_8 : in std_logic_vector( 16-1 downto 0 );
    in_9 : in std_logic_vector( 16-1 downto 0 );
    in_10 : in std_logic_vector( 16-1 downto 0 );
    in_11 : in std_logic_vector( 16-1 downto 0 );
    in_12 : in std_logic_vector( 16-1 downto 0 );
    in_13 : in std_logic_vector( 16-1 downto 0 );
    in_14 : in std_logic_vector( 16-1 downto 0 );
    in_15 : in std_logic_vector( 16-1 downto 0 );
    in_16 : in std_logic_vector( 16-1 downto 0 );
    out_1 : out std_logic_vector( 16-1 downto 0 );
    out_2 : out std_logic_vector( 16-1 downto 0 );
    out_3 : out std_logic_vector( 16-1 downto 0 );
    out_4 : out std_logic_vector( 16-1 downto 0 );
    out_5 : out std_logic_vector( 16-1 downto 0 );
    out_6 : out std_logic_vector( 16-1 downto 0 );
    out_7 : out std_logic_vector( 16-1 downto 0 );
    out_8 : out std_logic_vector( 16-1 downto 0 );
    out_9 : out std_logic_vector( 16-1 downto 0 );
    out_10 : out std_logic_vector( 16-1 downto 0 );
    out_11 : out std_logic_vector( 16-1 downto 0 );
    out_12 : out std_logic_vector( 16-1 downto 0 );
    out_13 : out std_logic_vector( 16-1 downto 0 );
    out_14 : out std_logic_vector( 16-1 downto 0 );
    out_15 : out std_logic_vector( 16-1 downto 0 );
    out_16 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_vector_reinterpret1;
architecture structural of psb3_0_vector_reinterpret1 is 
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 16-1 downto 0 );
begin
  out_1 <= reinterpret0_output_port_net;
  out_2 <= reinterpret1_output_port_net;
  out_3 <= reinterpret2_output_port_net;
  out_4 <= reinterpret3_output_port_net;
  out_5 <= reinterpret4_output_port_net;
  out_6 <= reinterpret5_output_port_net;
  out_7 <= reinterpret6_output_port_net;
  out_8 <= reinterpret7_output_port_net;
  out_9 <= reinterpret8_output_port_net;
  out_10 <= reinterpret9_output_port_net;
  out_11 <= reinterpret10_output_port_net;
  out_12 <= reinterpret11_output_port_net;
  out_13 <= reinterpret12_output_port_net;
  out_14 <= reinterpret13_output_port_net;
  out_15 <= reinterpret14_output_port_net;
  out_16 <= reinterpret15_output_port_net;
  slice0_y_net <= in_1;
  slice1_y_net <= in_2;
  slice2_y_net <= in_3;
  slice3_y_net <= in_4;
  slice4_y_net <= in_5;
  slice5_y_net <= in_6;
  slice6_y_net <= in_7;
  slice7_y_net <= in_8;
  slice8_y_net <= in_9;
  slice9_y_net <= in_10;
  slice10_y_net <= in_11;
  slice11_y_net <= in_12;
  slice12_y_net <= in_13;
  slice13_y_net <= in_14;
  slice14_y_net <= in_15;
  slice15_y_net <= in_16;
  reinterpret0 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice0_y_net,
    output_port => reinterpret0_output_port_net
  );
  reinterpret1 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice1_y_net,
    output_port => reinterpret1_output_port_net
  );
  reinterpret2 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice2_y_net,
    output_port => reinterpret2_output_port_net
  );
  reinterpret3 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice3_y_net,
    output_port => reinterpret3_output_port_net
  );
  reinterpret4 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice4_y_net,
    output_port => reinterpret4_output_port_net
  );
  reinterpret5 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice5_y_net,
    output_port => reinterpret5_output_port_net
  );
  reinterpret6 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice6_y_net,
    output_port => reinterpret6_output_port_net
  );
  reinterpret7 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice7_y_net,
    output_port => reinterpret7_output_port_net
  );
  reinterpret8 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice8_y_net,
    output_port => reinterpret8_output_port_net
  );
  reinterpret9 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice9_y_net,
    output_port => reinterpret9_output_port_net
  );
  reinterpret10 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice10_y_net,
    output_port => reinterpret10_output_port_net
  );
  reinterpret11 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice11_y_net,
    output_port => reinterpret11_output_port_net
  );
  reinterpret12 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice12_y_net,
    output_port => reinterpret12_output_port_net
  );
  reinterpret13 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice13_y_net,
    output_port => reinterpret13_output_port_net
  );
  reinterpret14 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice14_y_net,
    output_port => reinterpret14_output_port_net
  );
  reinterpret15 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice15_y_net,
    output_port => reinterpret15_output_port_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Vector Reinterpret10
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_reinterpret10 is
  port (
    in_1 : in std_logic_vector( 16-1 downto 0 );
    in_2 : in std_logic_vector( 16-1 downto 0 );
    in_3 : in std_logic_vector( 16-1 downto 0 );
    in_4 : in std_logic_vector( 16-1 downto 0 );
    in_5 : in std_logic_vector( 16-1 downto 0 );
    in_6 : in std_logic_vector( 16-1 downto 0 );
    in_7 : in std_logic_vector( 16-1 downto 0 );
    in_8 : in std_logic_vector( 16-1 downto 0 );
    in_9 : in std_logic_vector( 16-1 downto 0 );
    in_10 : in std_logic_vector( 16-1 downto 0 );
    in_11 : in std_logic_vector( 16-1 downto 0 );
    in_12 : in std_logic_vector( 16-1 downto 0 );
    in_13 : in std_logic_vector( 16-1 downto 0 );
    in_14 : in std_logic_vector( 16-1 downto 0 );
    in_15 : in std_logic_vector( 16-1 downto 0 );
    in_16 : in std_logic_vector( 16-1 downto 0 );
    out_1 : out std_logic_vector( 16-1 downto 0 );
    out_2 : out std_logic_vector( 16-1 downto 0 );
    out_3 : out std_logic_vector( 16-1 downto 0 );
    out_4 : out std_logic_vector( 16-1 downto 0 );
    out_5 : out std_logic_vector( 16-1 downto 0 );
    out_6 : out std_logic_vector( 16-1 downto 0 );
    out_7 : out std_logic_vector( 16-1 downto 0 );
    out_8 : out std_logic_vector( 16-1 downto 0 );
    out_9 : out std_logic_vector( 16-1 downto 0 );
    out_10 : out std_logic_vector( 16-1 downto 0 );
    out_11 : out std_logic_vector( 16-1 downto 0 );
    out_12 : out std_logic_vector( 16-1 downto 0 );
    out_13 : out std_logic_vector( 16-1 downto 0 );
    out_14 : out std_logic_vector( 16-1 downto 0 );
    out_15 : out std_logic_vector( 16-1 downto 0 );
    out_16 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_vector_reinterpret10;
architecture structural of psb3_0_vector_reinterpret10 is 
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
begin
  out_1 <= reinterpret0_output_port_net;
  out_2 <= reinterpret1_output_port_net;
  out_3 <= reinterpret2_output_port_net;
  out_4 <= reinterpret3_output_port_net;
  out_5 <= reinterpret4_output_port_net;
  out_6 <= reinterpret5_output_port_net;
  out_7 <= reinterpret6_output_port_net;
  out_8 <= reinterpret7_output_port_net;
  out_9 <= reinterpret8_output_port_net;
  out_10 <= reinterpret9_output_port_net;
  out_11 <= reinterpret10_output_port_net;
  out_12 <= reinterpret11_output_port_net;
  out_13 <= reinterpret12_output_port_net;
  out_14 <= reinterpret13_output_port_net;
  out_15 <= reinterpret14_output_port_net;
  out_16 <= reinterpret15_output_port_net;
  slice0_y_net <= in_1;
  slice1_y_net <= in_2;
  slice2_y_net <= in_3;
  slice3_y_net <= in_4;
  slice4_y_net <= in_5;
  slice5_y_net <= in_6;
  slice6_y_net <= in_7;
  slice7_y_net <= in_8;
  slice8_y_net <= in_9;
  slice9_y_net <= in_10;
  slice10_y_net <= in_11;
  slice11_y_net <= in_12;
  slice12_y_net <= in_13;
  slice13_y_net <= in_14;
  slice14_y_net <= in_15;
  slice15_y_net <= in_16;
  reinterpret0 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice0_y_net,
    output_port => reinterpret0_output_port_net
  );
  reinterpret1 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice1_y_net,
    output_port => reinterpret1_output_port_net
  );
  reinterpret2 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice2_y_net,
    output_port => reinterpret2_output_port_net
  );
  reinterpret3 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice3_y_net,
    output_port => reinterpret3_output_port_net
  );
  reinterpret4 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice4_y_net,
    output_port => reinterpret4_output_port_net
  );
  reinterpret5 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice5_y_net,
    output_port => reinterpret5_output_port_net
  );
  reinterpret6 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice6_y_net,
    output_port => reinterpret6_output_port_net
  );
  reinterpret7 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice7_y_net,
    output_port => reinterpret7_output_port_net
  );
  reinterpret8 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice8_y_net,
    output_port => reinterpret8_output_port_net
  );
  reinterpret9 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice9_y_net,
    output_port => reinterpret9_output_port_net
  );
  reinterpret10 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice10_y_net,
    output_port => reinterpret10_output_port_net
  );
  reinterpret11 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice11_y_net,
    output_port => reinterpret11_output_port_net
  );
  reinterpret12 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice12_y_net,
    output_port => reinterpret12_output_port_net
  );
  reinterpret13 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice13_y_net,
    output_port => reinterpret13_output_port_net
  );
  reinterpret14 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice14_y_net,
    output_port => reinterpret14_output_port_net
  );
  reinterpret15 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice15_y_net,
    output_port => reinterpret15_output_port_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Vector Reinterpret11
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_reinterpret11 is
  port (
    in_1 : in std_logic_vector( 16-1 downto 0 );
    in_2 : in std_logic_vector( 16-1 downto 0 );
    in_3 : in std_logic_vector( 16-1 downto 0 );
    in_4 : in std_logic_vector( 16-1 downto 0 );
    in_5 : in std_logic_vector( 16-1 downto 0 );
    in_6 : in std_logic_vector( 16-1 downto 0 );
    in_7 : in std_logic_vector( 16-1 downto 0 );
    in_8 : in std_logic_vector( 16-1 downto 0 );
    in_9 : in std_logic_vector( 16-1 downto 0 );
    in_10 : in std_logic_vector( 16-1 downto 0 );
    in_11 : in std_logic_vector( 16-1 downto 0 );
    in_12 : in std_logic_vector( 16-1 downto 0 );
    in_13 : in std_logic_vector( 16-1 downto 0 );
    in_14 : in std_logic_vector( 16-1 downto 0 );
    in_15 : in std_logic_vector( 16-1 downto 0 );
    in_16 : in std_logic_vector( 16-1 downto 0 );
    out_1 : out std_logic_vector( 16-1 downto 0 );
    out_2 : out std_logic_vector( 16-1 downto 0 );
    out_3 : out std_logic_vector( 16-1 downto 0 );
    out_4 : out std_logic_vector( 16-1 downto 0 );
    out_5 : out std_logic_vector( 16-1 downto 0 );
    out_6 : out std_logic_vector( 16-1 downto 0 );
    out_7 : out std_logic_vector( 16-1 downto 0 );
    out_8 : out std_logic_vector( 16-1 downto 0 );
    out_9 : out std_logic_vector( 16-1 downto 0 );
    out_10 : out std_logic_vector( 16-1 downto 0 );
    out_11 : out std_logic_vector( 16-1 downto 0 );
    out_12 : out std_logic_vector( 16-1 downto 0 );
    out_13 : out std_logic_vector( 16-1 downto 0 );
    out_14 : out std_logic_vector( 16-1 downto 0 );
    out_15 : out std_logic_vector( 16-1 downto 0 );
    out_16 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_vector_reinterpret11;
architecture structural of psb3_0_vector_reinterpret11 is 
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 16-1 downto 0 );
begin
  out_1 <= reinterpret0_output_port_net;
  out_2 <= reinterpret1_output_port_net;
  out_3 <= reinterpret2_output_port_net;
  out_4 <= reinterpret3_output_port_net;
  out_5 <= reinterpret4_output_port_net;
  out_6 <= reinterpret5_output_port_net;
  out_7 <= reinterpret6_output_port_net;
  out_8 <= reinterpret7_output_port_net;
  out_9 <= reinterpret8_output_port_net;
  out_10 <= reinterpret9_output_port_net;
  out_11 <= reinterpret10_output_port_net;
  out_12 <= reinterpret11_output_port_net;
  out_13 <= reinterpret12_output_port_net;
  out_14 <= reinterpret13_output_port_net;
  out_15 <= reinterpret14_output_port_net;
  out_16 <= reinterpret15_output_port_net;
  slice0_y_net <= in_1;
  slice1_y_net <= in_2;
  slice2_y_net <= in_3;
  slice3_y_net <= in_4;
  slice4_y_net <= in_5;
  slice5_y_net <= in_6;
  slice6_y_net <= in_7;
  slice7_y_net <= in_8;
  slice8_y_net <= in_9;
  slice9_y_net <= in_10;
  slice10_y_net <= in_11;
  slice11_y_net <= in_12;
  slice12_y_net <= in_13;
  slice13_y_net <= in_14;
  slice14_y_net <= in_15;
  slice15_y_net <= in_16;
  reinterpret0 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice0_y_net,
    output_port => reinterpret0_output_port_net
  );
  reinterpret1 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice1_y_net,
    output_port => reinterpret1_output_port_net
  );
  reinterpret2 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice2_y_net,
    output_port => reinterpret2_output_port_net
  );
  reinterpret3 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice3_y_net,
    output_port => reinterpret3_output_port_net
  );
  reinterpret4 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice4_y_net,
    output_port => reinterpret4_output_port_net
  );
  reinterpret5 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice5_y_net,
    output_port => reinterpret5_output_port_net
  );
  reinterpret6 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice6_y_net,
    output_port => reinterpret6_output_port_net
  );
  reinterpret7 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice7_y_net,
    output_port => reinterpret7_output_port_net
  );
  reinterpret8 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice8_y_net,
    output_port => reinterpret8_output_port_net
  );
  reinterpret9 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice9_y_net,
    output_port => reinterpret9_output_port_net
  );
  reinterpret10 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice10_y_net,
    output_port => reinterpret10_output_port_net
  );
  reinterpret11 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice11_y_net,
    output_port => reinterpret11_output_port_net
  );
  reinterpret12 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice12_y_net,
    output_port => reinterpret12_output_port_net
  );
  reinterpret13 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice13_y_net,
    output_port => reinterpret13_output_port_net
  );
  reinterpret14 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice14_y_net,
    output_port => reinterpret14_output_port_net
  );
  reinterpret15 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice15_y_net,
    output_port => reinterpret15_output_port_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Vector Reinterpret12
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_reinterpret12 is
  port (
    in_1 : in std_logic_vector( 16-1 downto 0 );
    in_2 : in std_logic_vector( 16-1 downto 0 );
    in_3 : in std_logic_vector( 16-1 downto 0 );
    in_4 : in std_logic_vector( 16-1 downto 0 );
    in_5 : in std_logic_vector( 16-1 downto 0 );
    in_6 : in std_logic_vector( 16-1 downto 0 );
    in_7 : in std_logic_vector( 16-1 downto 0 );
    in_8 : in std_logic_vector( 16-1 downto 0 );
    in_9 : in std_logic_vector( 16-1 downto 0 );
    in_10 : in std_logic_vector( 16-1 downto 0 );
    in_11 : in std_logic_vector( 16-1 downto 0 );
    in_12 : in std_logic_vector( 16-1 downto 0 );
    in_13 : in std_logic_vector( 16-1 downto 0 );
    in_14 : in std_logic_vector( 16-1 downto 0 );
    in_15 : in std_logic_vector( 16-1 downto 0 );
    in_16 : in std_logic_vector( 16-1 downto 0 );
    out_1 : out std_logic_vector( 16-1 downto 0 );
    out_2 : out std_logic_vector( 16-1 downto 0 );
    out_3 : out std_logic_vector( 16-1 downto 0 );
    out_4 : out std_logic_vector( 16-1 downto 0 );
    out_5 : out std_logic_vector( 16-1 downto 0 );
    out_6 : out std_logic_vector( 16-1 downto 0 );
    out_7 : out std_logic_vector( 16-1 downto 0 );
    out_8 : out std_logic_vector( 16-1 downto 0 );
    out_9 : out std_logic_vector( 16-1 downto 0 );
    out_10 : out std_logic_vector( 16-1 downto 0 );
    out_11 : out std_logic_vector( 16-1 downto 0 );
    out_12 : out std_logic_vector( 16-1 downto 0 );
    out_13 : out std_logic_vector( 16-1 downto 0 );
    out_14 : out std_logic_vector( 16-1 downto 0 );
    out_15 : out std_logic_vector( 16-1 downto 0 );
    out_16 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_vector_reinterpret12;
architecture structural of psb3_0_vector_reinterpret12 is 
  signal addsub5_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub6_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub7_s_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub8_s_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub9_s_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub0_s_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub3_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub12_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub14_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub10_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub15_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub13_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub11_s_net : std_logic_vector( 16-1 downto 0 );
begin
  out_1 <= reinterpret0_output_port_net;
  out_2 <= reinterpret1_output_port_net;
  out_3 <= reinterpret2_output_port_net;
  out_4 <= reinterpret3_output_port_net;
  out_5 <= reinterpret4_output_port_net;
  out_6 <= reinterpret5_output_port_net;
  out_7 <= reinterpret6_output_port_net;
  out_8 <= reinterpret7_output_port_net;
  out_9 <= reinterpret8_output_port_net;
  out_10 <= reinterpret9_output_port_net;
  out_11 <= reinterpret10_output_port_net;
  out_12 <= reinterpret11_output_port_net;
  out_13 <= reinterpret12_output_port_net;
  out_14 <= reinterpret13_output_port_net;
  out_15 <= reinterpret14_output_port_net;
  out_16 <= reinterpret15_output_port_net;
  addsub0_s_net <= in_1;
  addsub1_s_net <= in_2;
  addsub2_s_net <= in_3;
  addsub3_s_net <= in_4;
  addsub4_s_net <= in_5;
  addsub5_s_net <= in_6;
  addsub6_s_net <= in_7;
  addsub7_s_net <= in_8;
  addsub8_s_net <= in_9;
  addsub9_s_net <= in_10;
  addsub10_s_net <= in_11;
  addsub11_s_net <= in_12;
  addsub12_s_net <= in_13;
  addsub13_s_net <= in_14;
  addsub14_s_net <= in_15;
  addsub15_s_net <= in_16;
  reinterpret0 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub0_s_net,
    output_port => reinterpret0_output_port_net
  );
  reinterpret1 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub1_s_net,
    output_port => reinterpret1_output_port_net
  );
  reinterpret2 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub2_s_net,
    output_port => reinterpret2_output_port_net
  );
  reinterpret3 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub3_s_net,
    output_port => reinterpret3_output_port_net
  );
  reinterpret4 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub4_s_net,
    output_port => reinterpret4_output_port_net
  );
  reinterpret5 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub5_s_net,
    output_port => reinterpret5_output_port_net
  );
  reinterpret6 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub6_s_net,
    output_port => reinterpret6_output_port_net
  );
  reinterpret7 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub7_s_net,
    output_port => reinterpret7_output_port_net
  );
  reinterpret8 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub8_s_net,
    output_port => reinterpret8_output_port_net
  );
  reinterpret9 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub9_s_net,
    output_port => reinterpret9_output_port_net
  );
  reinterpret10 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub10_s_net,
    output_port => reinterpret10_output_port_net
  );
  reinterpret11 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub11_s_net,
    output_port => reinterpret11_output_port_net
  );
  reinterpret12 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub12_s_net,
    output_port => reinterpret12_output_port_net
  );
  reinterpret13 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub13_s_net,
    output_port => reinterpret13_output_port_net
  );
  reinterpret14 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub14_s_net,
    output_port => reinterpret14_output_port_net
  );
  reinterpret15 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub15_s_net,
    output_port => reinterpret15_output_port_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Vector Reinterpret13
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_reinterpret13 is
  port (
    in_1 : in std_logic_vector( 16-1 downto 0 );
    in_2 : in std_logic_vector( 16-1 downto 0 );
    in_3 : in std_logic_vector( 16-1 downto 0 );
    in_4 : in std_logic_vector( 16-1 downto 0 );
    in_5 : in std_logic_vector( 16-1 downto 0 );
    in_6 : in std_logic_vector( 16-1 downto 0 );
    in_7 : in std_logic_vector( 16-1 downto 0 );
    in_8 : in std_logic_vector( 16-1 downto 0 );
    in_9 : in std_logic_vector( 16-1 downto 0 );
    in_10 : in std_logic_vector( 16-1 downto 0 );
    in_11 : in std_logic_vector( 16-1 downto 0 );
    in_12 : in std_logic_vector( 16-1 downto 0 );
    in_13 : in std_logic_vector( 16-1 downto 0 );
    in_14 : in std_logic_vector( 16-1 downto 0 );
    in_15 : in std_logic_vector( 16-1 downto 0 );
    in_16 : in std_logic_vector( 16-1 downto 0 );
    out_1 : out std_logic_vector( 16-1 downto 0 );
    out_2 : out std_logic_vector( 16-1 downto 0 );
    out_3 : out std_logic_vector( 16-1 downto 0 );
    out_4 : out std_logic_vector( 16-1 downto 0 );
    out_5 : out std_logic_vector( 16-1 downto 0 );
    out_6 : out std_logic_vector( 16-1 downto 0 );
    out_7 : out std_logic_vector( 16-1 downto 0 );
    out_8 : out std_logic_vector( 16-1 downto 0 );
    out_9 : out std_logic_vector( 16-1 downto 0 );
    out_10 : out std_logic_vector( 16-1 downto 0 );
    out_11 : out std_logic_vector( 16-1 downto 0 );
    out_12 : out std_logic_vector( 16-1 downto 0 );
    out_13 : out std_logic_vector( 16-1 downto 0 );
    out_14 : out std_logic_vector( 16-1 downto 0 );
    out_15 : out std_logic_vector( 16-1 downto 0 );
    out_16 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_vector_reinterpret13;
architecture structural of psb3_0_vector_reinterpret13 is 
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub0_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub12_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub13_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub15_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub10_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub14_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub3_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub6_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub8_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub7_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub11_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub5_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub9_s_net : std_logic_vector( 16-1 downto 0 );
begin
  out_1 <= reinterpret0_output_port_net;
  out_2 <= reinterpret1_output_port_net;
  out_3 <= reinterpret2_output_port_net;
  out_4 <= reinterpret3_output_port_net;
  out_5 <= reinterpret4_output_port_net;
  out_6 <= reinterpret5_output_port_net;
  out_7 <= reinterpret6_output_port_net;
  out_8 <= reinterpret7_output_port_net;
  out_9 <= reinterpret8_output_port_net;
  out_10 <= reinterpret9_output_port_net;
  out_11 <= reinterpret10_output_port_net;
  out_12 <= reinterpret11_output_port_net;
  out_13 <= reinterpret12_output_port_net;
  out_14 <= reinterpret13_output_port_net;
  out_15 <= reinterpret14_output_port_net;
  out_16 <= reinterpret15_output_port_net;
  addsub0_s_net <= in_1;
  addsub1_s_net <= in_2;
  addsub2_s_net <= in_3;
  addsub3_s_net <= in_4;
  addsub4_s_net <= in_5;
  addsub5_s_net <= in_6;
  addsub6_s_net <= in_7;
  addsub7_s_net <= in_8;
  addsub8_s_net <= in_9;
  addsub9_s_net <= in_10;
  addsub10_s_net <= in_11;
  addsub11_s_net <= in_12;
  addsub12_s_net <= in_13;
  addsub13_s_net <= in_14;
  addsub14_s_net <= in_15;
  addsub15_s_net <= in_16;
  reinterpret0 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub0_s_net,
    output_port => reinterpret0_output_port_net
  );
  reinterpret1 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub1_s_net,
    output_port => reinterpret1_output_port_net
  );
  reinterpret2 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub2_s_net,
    output_port => reinterpret2_output_port_net
  );
  reinterpret3 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub3_s_net,
    output_port => reinterpret3_output_port_net
  );
  reinterpret4 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub4_s_net,
    output_port => reinterpret4_output_port_net
  );
  reinterpret5 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub5_s_net,
    output_port => reinterpret5_output_port_net
  );
  reinterpret6 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub6_s_net,
    output_port => reinterpret6_output_port_net
  );
  reinterpret7 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub7_s_net,
    output_port => reinterpret7_output_port_net
  );
  reinterpret8 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub8_s_net,
    output_port => reinterpret8_output_port_net
  );
  reinterpret9 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub9_s_net,
    output_port => reinterpret9_output_port_net
  );
  reinterpret10 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub10_s_net,
    output_port => reinterpret10_output_port_net
  );
  reinterpret11 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub11_s_net,
    output_port => reinterpret11_output_port_net
  );
  reinterpret12 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub12_s_net,
    output_port => reinterpret12_output_port_net
  );
  reinterpret13 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub13_s_net,
    output_port => reinterpret13_output_port_net
  );
  reinterpret14 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub14_s_net,
    output_port => reinterpret14_output_port_net
  );
  reinterpret15 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub15_s_net,
    output_port => reinterpret15_output_port_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Vector Reinterpret14
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_reinterpret14 is
  port (
    in_1 : in std_logic_vector( 16-1 downto 0 );
    in_2 : in std_logic_vector( 16-1 downto 0 );
    in_3 : in std_logic_vector( 16-1 downto 0 );
    in_4 : in std_logic_vector( 16-1 downto 0 );
    in_5 : in std_logic_vector( 16-1 downto 0 );
    in_6 : in std_logic_vector( 16-1 downto 0 );
    in_7 : in std_logic_vector( 16-1 downto 0 );
    in_8 : in std_logic_vector( 16-1 downto 0 );
    in_9 : in std_logic_vector( 16-1 downto 0 );
    in_10 : in std_logic_vector( 16-1 downto 0 );
    in_11 : in std_logic_vector( 16-1 downto 0 );
    in_12 : in std_logic_vector( 16-1 downto 0 );
    in_13 : in std_logic_vector( 16-1 downto 0 );
    in_14 : in std_logic_vector( 16-1 downto 0 );
    in_15 : in std_logic_vector( 16-1 downto 0 );
    in_16 : in std_logic_vector( 16-1 downto 0 );
    out_1 : out std_logic_vector( 16-1 downto 0 );
    out_2 : out std_logic_vector( 16-1 downto 0 );
    out_3 : out std_logic_vector( 16-1 downto 0 );
    out_4 : out std_logic_vector( 16-1 downto 0 );
    out_5 : out std_logic_vector( 16-1 downto 0 );
    out_6 : out std_logic_vector( 16-1 downto 0 );
    out_7 : out std_logic_vector( 16-1 downto 0 );
    out_8 : out std_logic_vector( 16-1 downto 0 );
    out_9 : out std_logic_vector( 16-1 downto 0 );
    out_10 : out std_logic_vector( 16-1 downto 0 );
    out_11 : out std_logic_vector( 16-1 downto 0 );
    out_12 : out std_logic_vector( 16-1 downto 0 );
    out_13 : out std_logic_vector( 16-1 downto 0 );
    out_14 : out std_logic_vector( 16-1 downto 0 );
    out_15 : out std_logic_vector( 16-1 downto 0 );
    out_16 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_vector_reinterpret14;
architecture structural of psb3_0_vector_reinterpret14 is 
  signal slice7_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
begin
  out_1 <= reinterpret0_output_port_net;
  out_2 <= reinterpret1_output_port_net;
  out_3 <= reinterpret2_output_port_net;
  out_4 <= reinterpret3_output_port_net;
  out_5 <= reinterpret4_output_port_net;
  out_6 <= reinterpret5_output_port_net;
  out_7 <= reinterpret6_output_port_net;
  out_8 <= reinterpret7_output_port_net;
  out_9 <= reinterpret8_output_port_net;
  out_10 <= reinterpret9_output_port_net;
  out_11 <= reinterpret10_output_port_net;
  out_12 <= reinterpret11_output_port_net;
  out_13 <= reinterpret12_output_port_net;
  out_14 <= reinterpret13_output_port_net;
  out_15 <= reinterpret14_output_port_net;
  out_16 <= reinterpret15_output_port_net;
  slice0_y_net <= in_1;
  slice1_y_net <= in_2;
  slice2_y_net <= in_3;
  slice3_y_net <= in_4;
  slice4_y_net <= in_5;
  slice5_y_net <= in_6;
  slice6_y_net <= in_7;
  slice7_y_net <= in_8;
  slice8_y_net <= in_9;
  slice9_y_net <= in_10;
  slice10_y_net <= in_11;
  slice11_y_net <= in_12;
  slice12_y_net <= in_13;
  slice13_y_net <= in_14;
  slice14_y_net <= in_15;
  slice15_y_net <= in_16;
  reinterpret0 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice0_y_net,
    output_port => reinterpret0_output_port_net
  );
  reinterpret1 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice1_y_net,
    output_port => reinterpret1_output_port_net
  );
  reinterpret2 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice2_y_net,
    output_port => reinterpret2_output_port_net
  );
  reinterpret3 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice3_y_net,
    output_port => reinterpret3_output_port_net
  );
  reinterpret4 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice4_y_net,
    output_port => reinterpret4_output_port_net
  );
  reinterpret5 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice5_y_net,
    output_port => reinterpret5_output_port_net
  );
  reinterpret6 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice6_y_net,
    output_port => reinterpret6_output_port_net
  );
  reinterpret7 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice7_y_net,
    output_port => reinterpret7_output_port_net
  );
  reinterpret8 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice8_y_net,
    output_port => reinterpret8_output_port_net
  );
  reinterpret9 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice9_y_net,
    output_port => reinterpret9_output_port_net
  );
  reinterpret10 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice10_y_net,
    output_port => reinterpret10_output_port_net
  );
  reinterpret11 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice11_y_net,
    output_port => reinterpret11_output_port_net
  );
  reinterpret12 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice12_y_net,
    output_port => reinterpret12_output_port_net
  );
  reinterpret13 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice13_y_net,
    output_port => reinterpret13_output_port_net
  );
  reinterpret14 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice14_y_net,
    output_port => reinterpret14_output_port_net
  );
  reinterpret15 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice15_y_net,
    output_port => reinterpret15_output_port_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Vector Reinterpret15
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_reinterpret15 is
  port (
    in_1 : in std_logic_vector( 16-1 downto 0 );
    in_2 : in std_logic_vector( 16-1 downto 0 );
    in_3 : in std_logic_vector( 16-1 downto 0 );
    in_4 : in std_logic_vector( 16-1 downto 0 );
    in_5 : in std_logic_vector( 16-1 downto 0 );
    in_6 : in std_logic_vector( 16-1 downto 0 );
    in_7 : in std_logic_vector( 16-1 downto 0 );
    in_8 : in std_logic_vector( 16-1 downto 0 );
    in_9 : in std_logic_vector( 16-1 downto 0 );
    in_10 : in std_logic_vector( 16-1 downto 0 );
    in_11 : in std_logic_vector( 16-1 downto 0 );
    in_12 : in std_logic_vector( 16-1 downto 0 );
    in_13 : in std_logic_vector( 16-1 downto 0 );
    in_14 : in std_logic_vector( 16-1 downto 0 );
    in_15 : in std_logic_vector( 16-1 downto 0 );
    in_16 : in std_logic_vector( 16-1 downto 0 );
    out_1 : out std_logic_vector( 16-1 downto 0 );
    out_2 : out std_logic_vector( 16-1 downto 0 );
    out_3 : out std_logic_vector( 16-1 downto 0 );
    out_4 : out std_logic_vector( 16-1 downto 0 );
    out_5 : out std_logic_vector( 16-1 downto 0 );
    out_6 : out std_logic_vector( 16-1 downto 0 );
    out_7 : out std_logic_vector( 16-1 downto 0 );
    out_8 : out std_logic_vector( 16-1 downto 0 );
    out_9 : out std_logic_vector( 16-1 downto 0 );
    out_10 : out std_logic_vector( 16-1 downto 0 );
    out_11 : out std_logic_vector( 16-1 downto 0 );
    out_12 : out std_logic_vector( 16-1 downto 0 );
    out_13 : out std_logic_vector( 16-1 downto 0 );
    out_14 : out std_logic_vector( 16-1 downto 0 );
    out_15 : out std_logic_vector( 16-1 downto 0 );
    out_16 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_vector_reinterpret15;
architecture structural of psb3_0_vector_reinterpret15 is 
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub12_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub5_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub13_s_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub14_s_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub3_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub6_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub7_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub8_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub9_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub11_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub10_s_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub0_s_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub15_s_net : std_logic_vector( 16-1 downto 0 );
begin
  out_1 <= reinterpret0_output_port_net;
  out_2 <= reinterpret1_output_port_net;
  out_3 <= reinterpret2_output_port_net;
  out_4 <= reinterpret3_output_port_net;
  out_5 <= reinterpret4_output_port_net;
  out_6 <= reinterpret5_output_port_net;
  out_7 <= reinterpret6_output_port_net;
  out_8 <= reinterpret7_output_port_net;
  out_9 <= reinterpret8_output_port_net;
  out_10 <= reinterpret9_output_port_net;
  out_11 <= reinterpret10_output_port_net;
  out_12 <= reinterpret11_output_port_net;
  out_13 <= reinterpret12_output_port_net;
  out_14 <= reinterpret13_output_port_net;
  out_15 <= reinterpret14_output_port_net;
  out_16 <= reinterpret15_output_port_net;
  addsub0_s_net <= in_1;
  addsub1_s_net <= in_2;
  addsub2_s_net <= in_3;
  addsub3_s_net <= in_4;
  addsub4_s_net <= in_5;
  addsub5_s_net <= in_6;
  addsub6_s_net <= in_7;
  addsub7_s_net <= in_8;
  addsub8_s_net <= in_9;
  addsub9_s_net <= in_10;
  addsub10_s_net <= in_11;
  addsub11_s_net <= in_12;
  addsub12_s_net <= in_13;
  addsub13_s_net <= in_14;
  addsub14_s_net <= in_15;
  addsub15_s_net <= in_16;
  reinterpret0 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub0_s_net,
    output_port => reinterpret0_output_port_net
  );
  reinterpret1 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub1_s_net,
    output_port => reinterpret1_output_port_net
  );
  reinterpret2 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub2_s_net,
    output_port => reinterpret2_output_port_net
  );
  reinterpret3 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub3_s_net,
    output_port => reinterpret3_output_port_net
  );
  reinterpret4 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub4_s_net,
    output_port => reinterpret4_output_port_net
  );
  reinterpret5 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub5_s_net,
    output_port => reinterpret5_output_port_net
  );
  reinterpret6 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub6_s_net,
    output_port => reinterpret6_output_port_net
  );
  reinterpret7 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub7_s_net,
    output_port => reinterpret7_output_port_net
  );
  reinterpret8 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub8_s_net,
    output_port => reinterpret8_output_port_net
  );
  reinterpret9 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub9_s_net,
    output_port => reinterpret9_output_port_net
  );
  reinterpret10 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub10_s_net,
    output_port => reinterpret10_output_port_net
  );
  reinterpret11 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub11_s_net,
    output_port => reinterpret11_output_port_net
  );
  reinterpret12 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub12_s_net,
    output_port => reinterpret12_output_port_net
  );
  reinterpret13 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub13_s_net,
    output_port => reinterpret13_output_port_net
  );
  reinterpret14 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub14_s_net,
    output_port => reinterpret14_output_port_net
  );
  reinterpret15 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub15_s_net,
    output_port => reinterpret15_output_port_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Vector Reinterpret16
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_reinterpret16 is
  port (
    in_1 : in std_logic_vector( 16-1 downto 0 );
    in_2 : in std_logic_vector( 16-1 downto 0 );
    in_3 : in std_logic_vector( 16-1 downto 0 );
    in_4 : in std_logic_vector( 16-1 downto 0 );
    in_5 : in std_logic_vector( 16-1 downto 0 );
    in_6 : in std_logic_vector( 16-1 downto 0 );
    in_7 : in std_logic_vector( 16-1 downto 0 );
    in_8 : in std_logic_vector( 16-1 downto 0 );
    in_9 : in std_logic_vector( 16-1 downto 0 );
    in_10 : in std_logic_vector( 16-1 downto 0 );
    in_11 : in std_logic_vector( 16-1 downto 0 );
    in_12 : in std_logic_vector( 16-1 downto 0 );
    in_13 : in std_logic_vector( 16-1 downto 0 );
    in_14 : in std_logic_vector( 16-1 downto 0 );
    in_15 : in std_logic_vector( 16-1 downto 0 );
    in_16 : in std_logic_vector( 16-1 downto 0 );
    out_1 : out std_logic_vector( 16-1 downto 0 );
    out_2 : out std_logic_vector( 16-1 downto 0 );
    out_3 : out std_logic_vector( 16-1 downto 0 );
    out_4 : out std_logic_vector( 16-1 downto 0 );
    out_5 : out std_logic_vector( 16-1 downto 0 );
    out_6 : out std_logic_vector( 16-1 downto 0 );
    out_7 : out std_logic_vector( 16-1 downto 0 );
    out_8 : out std_logic_vector( 16-1 downto 0 );
    out_9 : out std_logic_vector( 16-1 downto 0 );
    out_10 : out std_logic_vector( 16-1 downto 0 );
    out_11 : out std_logic_vector( 16-1 downto 0 );
    out_12 : out std_logic_vector( 16-1 downto 0 );
    out_13 : out std_logic_vector( 16-1 downto 0 );
    out_14 : out std_logic_vector( 16-1 downto 0 );
    out_15 : out std_logic_vector( 16-1 downto 0 );
    out_16 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_vector_reinterpret16;
architecture structural of psb3_0_vector_reinterpret16 is 
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub5_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub6_s_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub0_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub3_s_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub13_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub9_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub12_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub14_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub15_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub8_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub7_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub11_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub10_s_net : std_logic_vector( 16-1 downto 0 );
begin
  out_1 <= reinterpret0_output_port_net;
  out_2 <= reinterpret1_output_port_net;
  out_3 <= reinterpret2_output_port_net;
  out_4 <= reinterpret3_output_port_net;
  out_5 <= reinterpret4_output_port_net;
  out_6 <= reinterpret5_output_port_net;
  out_7 <= reinterpret6_output_port_net;
  out_8 <= reinterpret7_output_port_net;
  out_9 <= reinterpret8_output_port_net;
  out_10 <= reinterpret9_output_port_net;
  out_11 <= reinterpret10_output_port_net;
  out_12 <= reinterpret11_output_port_net;
  out_13 <= reinterpret12_output_port_net;
  out_14 <= reinterpret13_output_port_net;
  out_15 <= reinterpret14_output_port_net;
  out_16 <= reinterpret15_output_port_net;
  addsub0_s_net <= in_1;
  addsub1_s_net <= in_2;
  addsub2_s_net <= in_3;
  addsub3_s_net <= in_4;
  addsub4_s_net <= in_5;
  addsub5_s_net <= in_6;
  addsub6_s_net <= in_7;
  addsub7_s_net <= in_8;
  addsub8_s_net <= in_9;
  addsub9_s_net <= in_10;
  addsub10_s_net <= in_11;
  addsub11_s_net <= in_12;
  addsub12_s_net <= in_13;
  addsub13_s_net <= in_14;
  addsub14_s_net <= in_15;
  addsub15_s_net <= in_16;
  reinterpret0 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub0_s_net,
    output_port => reinterpret0_output_port_net
  );
  reinterpret1 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub1_s_net,
    output_port => reinterpret1_output_port_net
  );
  reinterpret2 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub2_s_net,
    output_port => reinterpret2_output_port_net
  );
  reinterpret3 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub3_s_net,
    output_port => reinterpret3_output_port_net
  );
  reinterpret4 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub4_s_net,
    output_port => reinterpret4_output_port_net
  );
  reinterpret5 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub5_s_net,
    output_port => reinterpret5_output_port_net
  );
  reinterpret6 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub6_s_net,
    output_port => reinterpret6_output_port_net
  );
  reinterpret7 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub7_s_net,
    output_port => reinterpret7_output_port_net
  );
  reinterpret8 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub8_s_net,
    output_port => reinterpret8_output_port_net
  );
  reinterpret9 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub9_s_net,
    output_port => reinterpret9_output_port_net
  );
  reinterpret10 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub10_s_net,
    output_port => reinterpret10_output_port_net
  );
  reinterpret11 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub11_s_net,
    output_port => reinterpret11_output_port_net
  );
  reinterpret12 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub12_s_net,
    output_port => reinterpret12_output_port_net
  );
  reinterpret13 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub13_s_net,
    output_port => reinterpret13_output_port_net
  );
  reinterpret14 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub14_s_net,
    output_port => reinterpret14_output_port_net
  );
  reinterpret15 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub15_s_net,
    output_port => reinterpret15_output_port_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Vector Reinterpret2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_reinterpret2 is
  port (
    in_1 : in std_logic_vector( 16-1 downto 0 );
    in_2 : in std_logic_vector( 16-1 downto 0 );
    in_3 : in std_logic_vector( 16-1 downto 0 );
    in_4 : in std_logic_vector( 16-1 downto 0 );
    in_5 : in std_logic_vector( 16-1 downto 0 );
    in_6 : in std_logic_vector( 16-1 downto 0 );
    in_7 : in std_logic_vector( 16-1 downto 0 );
    in_8 : in std_logic_vector( 16-1 downto 0 );
    in_9 : in std_logic_vector( 16-1 downto 0 );
    in_10 : in std_logic_vector( 16-1 downto 0 );
    in_11 : in std_logic_vector( 16-1 downto 0 );
    in_12 : in std_logic_vector( 16-1 downto 0 );
    in_13 : in std_logic_vector( 16-1 downto 0 );
    in_14 : in std_logic_vector( 16-1 downto 0 );
    in_15 : in std_logic_vector( 16-1 downto 0 );
    in_16 : in std_logic_vector( 16-1 downto 0 );
    out_1 : out std_logic_vector( 16-1 downto 0 );
    out_2 : out std_logic_vector( 16-1 downto 0 );
    out_3 : out std_logic_vector( 16-1 downto 0 );
    out_4 : out std_logic_vector( 16-1 downto 0 );
    out_5 : out std_logic_vector( 16-1 downto 0 );
    out_6 : out std_logic_vector( 16-1 downto 0 );
    out_7 : out std_logic_vector( 16-1 downto 0 );
    out_8 : out std_logic_vector( 16-1 downto 0 );
    out_9 : out std_logic_vector( 16-1 downto 0 );
    out_10 : out std_logic_vector( 16-1 downto 0 );
    out_11 : out std_logic_vector( 16-1 downto 0 );
    out_12 : out std_logic_vector( 16-1 downto 0 );
    out_13 : out std_logic_vector( 16-1 downto 0 );
    out_14 : out std_logic_vector( 16-1 downto 0 );
    out_15 : out std_logic_vector( 16-1 downto 0 );
    out_16 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_vector_reinterpret2;
architecture structural of psb3_0_vector_reinterpret2 is 
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 16-1 downto 0 );
begin
  out_1 <= reinterpret0_output_port_net;
  out_2 <= reinterpret1_output_port_net;
  out_3 <= reinterpret2_output_port_net;
  out_4 <= reinterpret3_output_port_net;
  out_5 <= reinterpret4_output_port_net;
  out_6 <= reinterpret5_output_port_net;
  out_7 <= reinterpret6_output_port_net;
  out_8 <= reinterpret7_output_port_net;
  out_9 <= reinterpret8_output_port_net;
  out_10 <= reinterpret9_output_port_net;
  out_11 <= reinterpret10_output_port_net;
  out_12 <= reinterpret11_output_port_net;
  out_13 <= reinterpret12_output_port_net;
  out_14 <= reinterpret13_output_port_net;
  out_15 <= reinterpret14_output_port_net;
  out_16 <= reinterpret15_output_port_net;
  slice0_y_net <= in_1;
  slice1_y_net <= in_2;
  slice2_y_net <= in_3;
  slice3_y_net <= in_4;
  slice4_y_net <= in_5;
  slice5_y_net <= in_6;
  slice6_y_net <= in_7;
  slice7_y_net <= in_8;
  slice8_y_net <= in_9;
  slice9_y_net <= in_10;
  slice10_y_net <= in_11;
  slice11_y_net <= in_12;
  slice12_y_net <= in_13;
  slice13_y_net <= in_14;
  slice14_y_net <= in_15;
  slice15_y_net <= in_16;
  reinterpret0 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice0_y_net,
    output_port => reinterpret0_output_port_net
  );
  reinterpret1 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice1_y_net,
    output_port => reinterpret1_output_port_net
  );
  reinterpret2 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice2_y_net,
    output_port => reinterpret2_output_port_net
  );
  reinterpret3 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice3_y_net,
    output_port => reinterpret3_output_port_net
  );
  reinterpret4 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice4_y_net,
    output_port => reinterpret4_output_port_net
  );
  reinterpret5 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice5_y_net,
    output_port => reinterpret5_output_port_net
  );
  reinterpret6 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice6_y_net,
    output_port => reinterpret6_output_port_net
  );
  reinterpret7 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice7_y_net,
    output_port => reinterpret7_output_port_net
  );
  reinterpret8 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice8_y_net,
    output_port => reinterpret8_output_port_net
  );
  reinterpret9 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice9_y_net,
    output_port => reinterpret9_output_port_net
  );
  reinterpret10 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice10_y_net,
    output_port => reinterpret10_output_port_net
  );
  reinterpret11 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice11_y_net,
    output_port => reinterpret11_output_port_net
  );
  reinterpret12 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice12_y_net,
    output_port => reinterpret12_output_port_net
  );
  reinterpret13 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice13_y_net,
    output_port => reinterpret13_output_port_net
  );
  reinterpret14 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice14_y_net,
    output_port => reinterpret14_output_port_net
  );
  reinterpret15 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice15_y_net,
    output_port => reinterpret15_output_port_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Vector Reinterpret3
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_reinterpret3 is
  port (
    in_1 : in std_logic_vector( 16-1 downto 0 );
    in_2 : in std_logic_vector( 16-1 downto 0 );
    in_3 : in std_logic_vector( 16-1 downto 0 );
    in_4 : in std_logic_vector( 16-1 downto 0 );
    in_5 : in std_logic_vector( 16-1 downto 0 );
    in_6 : in std_logic_vector( 16-1 downto 0 );
    in_7 : in std_logic_vector( 16-1 downto 0 );
    in_8 : in std_logic_vector( 16-1 downto 0 );
    in_9 : in std_logic_vector( 16-1 downto 0 );
    in_10 : in std_logic_vector( 16-1 downto 0 );
    in_11 : in std_logic_vector( 16-1 downto 0 );
    in_12 : in std_logic_vector( 16-1 downto 0 );
    in_13 : in std_logic_vector( 16-1 downto 0 );
    in_14 : in std_logic_vector( 16-1 downto 0 );
    in_15 : in std_logic_vector( 16-1 downto 0 );
    in_16 : in std_logic_vector( 16-1 downto 0 );
    out_1 : out std_logic_vector( 16-1 downto 0 );
    out_2 : out std_logic_vector( 16-1 downto 0 );
    out_3 : out std_logic_vector( 16-1 downto 0 );
    out_4 : out std_logic_vector( 16-1 downto 0 );
    out_5 : out std_logic_vector( 16-1 downto 0 );
    out_6 : out std_logic_vector( 16-1 downto 0 );
    out_7 : out std_logic_vector( 16-1 downto 0 );
    out_8 : out std_logic_vector( 16-1 downto 0 );
    out_9 : out std_logic_vector( 16-1 downto 0 );
    out_10 : out std_logic_vector( 16-1 downto 0 );
    out_11 : out std_logic_vector( 16-1 downto 0 );
    out_12 : out std_logic_vector( 16-1 downto 0 );
    out_13 : out std_logic_vector( 16-1 downto 0 );
    out_14 : out std_logic_vector( 16-1 downto 0 );
    out_15 : out std_logic_vector( 16-1 downto 0 );
    out_16 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_vector_reinterpret3;
architecture structural of psb3_0_vector_reinterpret3 is 
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
begin
  out_1 <= reinterpret0_output_port_net;
  out_2 <= reinterpret1_output_port_net;
  out_3 <= reinterpret2_output_port_net;
  out_4 <= reinterpret3_output_port_net;
  out_5 <= reinterpret4_output_port_net;
  out_6 <= reinterpret5_output_port_net;
  out_7 <= reinterpret6_output_port_net;
  out_8 <= reinterpret7_output_port_net;
  out_9 <= reinterpret8_output_port_net;
  out_10 <= reinterpret9_output_port_net;
  out_11 <= reinterpret10_output_port_net;
  out_12 <= reinterpret11_output_port_net;
  out_13 <= reinterpret12_output_port_net;
  out_14 <= reinterpret13_output_port_net;
  out_15 <= reinterpret14_output_port_net;
  out_16 <= reinterpret15_output_port_net;
  slice0_y_net <= in_1;
  slice1_y_net <= in_2;
  slice2_y_net <= in_3;
  slice3_y_net <= in_4;
  slice4_y_net <= in_5;
  slice5_y_net <= in_6;
  slice6_y_net <= in_7;
  slice7_y_net <= in_8;
  slice8_y_net <= in_9;
  slice9_y_net <= in_10;
  slice10_y_net <= in_11;
  slice11_y_net <= in_12;
  slice12_y_net <= in_13;
  slice13_y_net <= in_14;
  slice14_y_net <= in_15;
  slice15_y_net <= in_16;
  reinterpret0 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice0_y_net,
    output_port => reinterpret0_output_port_net
  );
  reinterpret1 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice1_y_net,
    output_port => reinterpret1_output_port_net
  );
  reinterpret2 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice2_y_net,
    output_port => reinterpret2_output_port_net
  );
  reinterpret3 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice3_y_net,
    output_port => reinterpret3_output_port_net
  );
  reinterpret4 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice4_y_net,
    output_port => reinterpret4_output_port_net
  );
  reinterpret5 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice5_y_net,
    output_port => reinterpret5_output_port_net
  );
  reinterpret6 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice6_y_net,
    output_port => reinterpret6_output_port_net
  );
  reinterpret7 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice7_y_net,
    output_port => reinterpret7_output_port_net
  );
  reinterpret8 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice8_y_net,
    output_port => reinterpret8_output_port_net
  );
  reinterpret9 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice9_y_net,
    output_port => reinterpret9_output_port_net
  );
  reinterpret10 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice10_y_net,
    output_port => reinterpret10_output_port_net
  );
  reinterpret11 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice11_y_net,
    output_port => reinterpret11_output_port_net
  );
  reinterpret12 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice12_y_net,
    output_port => reinterpret12_output_port_net
  );
  reinterpret13 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice13_y_net,
    output_port => reinterpret13_output_port_net
  );
  reinterpret14 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice14_y_net,
    output_port => reinterpret14_output_port_net
  );
  reinterpret15 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice15_y_net,
    output_port => reinterpret15_output_port_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Vector Reinterpret4
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_reinterpret4 is
  port (
    in_1 : in std_logic_vector( 16-1 downto 0 );
    in_2 : in std_logic_vector( 16-1 downto 0 );
    in_3 : in std_logic_vector( 16-1 downto 0 );
    in_4 : in std_logic_vector( 16-1 downto 0 );
    in_5 : in std_logic_vector( 16-1 downto 0 );
    in_6 : in std_logic_vector( 16-1 downto 0 );
    in_7 : in std_logic_vector( 16-1 downto 0 );
    in_8 : in std_logic_vector( 16-1 downto 0 );
    in_9 : in std_logic_vector( 16-1 downto 0 );
    in_10 : in std_logic_vector( 16-1 downto 0 );
    in_11 : in std_logic_vector( 16-1 downto 0 );
    in_12 : in std_logic_vector( 16-1 downto 0 );
    in_13 : in std_logic_vector( 16-1 downto 0 );
    in_14 : in std_logic_vector( 16-1 downto 0 );
    in_15 : in std_logic_vector( 16-1 downto 0 );
    in_16 : in std_logic_vector( 16-1 downto 0 );
    out_1 : out std_logic_vector( 16-1 downto 0 );
    out_2 : out std_logic_vector( 16-1 downto 0 );
    out_3 : out std_logic_vector( 16-1 downto 0 );
    out_4 : out std_logic_vector( 16-1 downto 0 );
    out_5 : out std_logic_vector( 16-1 downto 0 );
    out_6 : out std_logic_vector( 16-1 downto 0 );
    out_7 : out std_logic_vector( 16-1 downto 0 );
    out_8 : out std_logic_vector( 16-1 downto 0 );
    out_9 : out std_logic_vector( 16-1 downto 0 );
    out_10 : out std_logic_vector( 16-1 downto 0 );
    out_11 : out std_logic_vector( 16-1 downto 0 );
    out_12 : out std_logic_vector( 16-1 downto 0 );
    out_13 : out std_logic_vector( 16-1 downto 0 );
    out_14 : out std_logic_vector( 16-1 downto 0 );
    out_15 : out std_logic_vector( 16-1 downto 0 );
    out_16 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_vector_reinterpret4;
architecture structural of psb3_0_vector_reinterpret4 is 
  signal addsub11_s_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub12_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub10_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub7_s_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub8_s_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub3_s_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub5_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub6_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub0_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub9_s_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub15_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub13_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub14_s_net : std_logic_vector( 16-1 downto 0 );
begin
  out_1 <= reinterpret0_output_port_net;
  out_2 <= reinterpret1_output_port_net;
  out_3 <= reinterpret2_output_port_net;
  out_4 <= reinterpret3_output_port_net;
  out_5 <= reinterpret4_output_port_net;
  out_6 <= reinterpret5_output_port_net;
  out_7 <= reinterpret6_output_port_net;
  out_8 <= reinterpret7_output_port_net;
  out_9 <= reinterpret8_output_port_net;
  out_10 <= reinterpret9_output_port_net;
  out_11 <= reinterpret10_output_port_net;
  out_12 <= reinterpret11_output_port_net;
  out_13 <= reinterpret12_output_port_net;
  out_14 <= reinterpret13_output_port_net;
  out_15 <= reinterpret14_output_port_net;
  out_16 <= reinterpret15_output_port_net;
  addsub0_s_net <= in_1;
  addsub1_s_net <= in_2;
  addsub2_s_net <= in_3;
  addsub3_s_net <= in_4;
  addsub4_s_net <= in_5;
  addsub5_s_net <= in_6;
  addsub6_s_net <= in_7;
  addsub7_s_net <= in_8;
  addsub8_s_net <= in_9;
  addsub9_s_net <= in_10;
  addsub10_s_net <= in_11;
  addsub11_s_net <= in_12;
  addsub12_s_net <= in_13;
  addsub13_s_net <= in_14;
  addsub14_s_net <= in_15;
  addsub15_s_net <= in_16;
  reinterpret0 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub0_s_net,
    output_port => reinterpret0_output_port_net
  );
  reinterpret1 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub1_s_net,
    output_port => reinterpret1_output_port_net
  );
  reinterpret2 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub2_s_net,
    output_port => reinterpret2_output_port_net
  );
  reinterpret3 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub3_s_net,
    output_port => reinterpret3_output_port_net
  );
  reinterpret4 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub4_s_net,
    output_port => reinterpret4_output_port_net
  );
  reinterpret5 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub5_s_net,
    output_port => reinterpret5_output_port_net
  );
  reinterpret6 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub6_s_net,
    output_port => reinterpret6_output_port_net
  );
  reinterpret7 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub7_s_net,
    output_port => reinterpret7_output_port_net
  );
  reinterpret8 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub8_s_net,
    output_port => reinterpret8_output_port_net
  );
  reinterpret9 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub9_s_net,
    output_port => reinterpret9_output_port_net
  );
  reinterpret10 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub10_s_net,
    output_port => reinterpret10_output_port_net
  );
  reinterpret11 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub11_s_net,
    output_port => reinterpret11_output_port_net
  );
  reinterpret12 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub12_s_net,
    output_port => reinterpret12_output_port_net
  );
  reinterpret13 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub13_s_net,
    output_port => reinterpret13_output_port_net
  );
  reinterpret14 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub14_s_net,
    output_port => reinterpret14_output_port_net
  );
  reinterpret15 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub15_s_net,
    output_port => reinterpret15_output_port_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Vector Reinterpret5
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_reinterpret5 is
  port (
    in_1 : in std_logic_vector( 16-1 downto 0 );
    in_2 : in std_logic_vector( 16-1 downto 0 );
    in_3 : in std_logic_vector( 16-1 downto 0 );
    in_4 : in std_logic_vector( 16-1 downto 0 );
    in_5 : in std_logic_vector( 16-1 downto 0 );
    in_6 : in std_logic_vector( 16-1 downto 0 );
    in_7 : in std_logic_vector( 16-1 downto 0 );
    in_8 : in std_logic_vector( 16-1 downto 0 );
    in_9 : in std_logic_vector( 16-1 downto 0 );
    in_10 : in std_logic_vector( 16-1 downto 0 );
    in_11 : in std_logic_vector( 16-1 downto 0 );
    in_12 : in std_logic_vector( 16-1 downto 0 );
    in_13 : in std_logic_vector( 16-1 downto 0 );
    in_14 : in std_logic_vector( 16-1 downto 0 );
    in_15 : in std_logic_vector( 16-1 downto 0 );
    in_16 : in std_logic_vector( 16-1 downto 0 );
    out_1 : out std_logic_vector( 16-1 downto 0 );
    out_2 : out std_logic_vector( 16-1 downto 0 );
    out_3 : out std_logic_vector( 16-1 downto 0 );
    out_4 : out std_logic_vector( 16-1 downto 0 );
    out_5 : out std_logic_vector( 16-1 downto 0 );
    out_6 : out std_logic_vector( 16-1 downto 0 );
    out_7 : out std_logic_vector( 16-1 downto 0 );
    out_8 : out std_logic_vector( 16-1 downto 0 );
    out_9 : out std_logic_vector( 16-1 downto 0 );
    out_10 : out std_logic_vector( 16-1 downto 0 );
    out_11 : out std_logic_vector( 16-1 downto 0 );
    out_12 : out std_logic_vector( 16-1 downto 0 );
    out_13 : out std_logic_vector( 16-1 downto 0 );
    out_14 : out std_logic_vector( 16-1 downto 0 );
    out_15 : out std_logic_vector( 16-1 downto 0 );
    out_16 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_vector_reinterpret5;
architecture structural of psb3_0_vector_reinterpret5 is 
  signal addsub2_s_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub3_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub0_s_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub11_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub10_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub12_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub8_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub14_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub6_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub9_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub13_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub5_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub15_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub7_s_net : std_logic_vector( 16-1 downto 0 );
begin
  out_1 <= reinterpret0_output_port_net;
  out_2 <= reinterpret1_output_port_net;
  out_3 <= reinterpret2_output_port_net;
  out_4 <= reinterpret3_output_port_net;
  out_5 <= reinterpret4_output_port_net;
  out_6 <= reinterpret5_output_port_net;
  out_7 <= reinterpret6_output_port_net;
  out_8 <= reinterpret7_output_port_net;
  out_9 <= reinterpret8_output_port_net;
  out_10 <= reinterpret9_output_port_net;
  out_11 <= reinterpret10_output_port_net;
  out_12 <= reinterpret11_output_port_net;
  out_13 <= reinterpret12_output_port_net;
  out_14 <= reinterpret13_output_port_net;
  out_15 <= reinterpret14_output_port_net;
  out_16 <= reinterpret15_output_port_net;
  addsub0_s_net <= in_1;
  addsub1_s_net <= in_2;
  addsub2_s_net <= in_3;
  addsub3_s_net <= in_4;
  addsub4_s_net <= in_5;
  addsub5_s_net <= in_6;
  addsub6_s_net <= in_7;
  addsub7_s_net <= in_8;
  addsub8_s_net <= in_9;
  addsub9_s_net <= in_10;
  addsub10_s_net <= in_11;
  addsub11_s_net <= in_12;
  addsub12_s_net <= in_13;
  addsub13_s_net <= in_14;
  addsub14_s_net <= in_15;
  addsub15_s_net <= in_16;
  reinterpret0 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub0_s_net,
    output_port => reinterpret0_output_port_net
  );
  reinterpret1 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub1_s_net,
    output_port => reinterpret1_output_port_net
  );
  reinterpret2 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub2_s_net,
    output_port => reinterpret2_output_port_net
  );
  reinterpret3 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub3_s_net,
    output_port => reinterpret3_output_port_net
  );
  reinterpret4 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub4_s_net,
    output_port => reinterpret4_output_port_net
  );
  reinterpret5 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub5_s_net,
    output_port => reinterpret5_output_port_net
  );
  reinterpret6 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub6_s_net,
    output_port => reinterpret6_output_port_net
  );
  reinterpret7 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub7_s_net,
    output_port => reinterpret7_output_port_net
  );
  reinterpret8 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub8_s_net,
    output_port => reinterpret8_output_port_net
  );
  reinterpret9 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub9_s_net,
    output_port => reinterpret9_output_port_net
  );
  reinterpret10 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub10_s_net,
    output_port => reinterpret10_output_port_net
  );
  reinterpret11 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub11_s_net,
    output_port => reinterpret11_output_port_net
  );
  reinterpret12 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub12_s_net,
    output_port => reinterpret12_output_port_net
  );
  reinterpret13 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub13_s_net,
    output_port => reinterpret13_output_port_net
  );
  reinterpret14 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub14_s_net,
    output_port => reinterpret14_output_port_net
  );
  reinterpret15 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub15_s_net,
    output_port => reinterpret15_output_port_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Vector Reinterpret6
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_reinterpret6 is
  port (
    in_1 : in std_logic_vector( 16-1 downto 0 );
    in_2 : in std_logic_vector( 16-1 downto 0 );
    in_3 : in std_logic_vector( 16-1 downto 0 );
    in_4 : in std_logic_vector( 16-1 downto 0 );
    in_5 : in std_logic_vector( 16-1 downto 0 );
    in_6 : in std_logic_vector( 16-1 downto 0 );
    in_7 : in std_logic_vector( 16-1 downto 0 );
    in_8 : in std_logic_vector( 16-1 downto 0 );
    in_9 : in std_logic_vector( 16-1 downto 0 );
    in_10 : in std_logic_vector( 16-1 downto 0 );
    in_11 : in std_logic_vector( 16-1 downto 0 );
    in_12 : in std_logic_vector( 16-1 downto 0 );
    in_13 : in std_logic_vector( 16-1 downto 0 );
    in_14 : in std_logic_vector( 16-1 downto 0 );
    in_15 : in std_logic_vector( 16-1 downto 0 );
    in_16 : in std_logic_vector( 16-1 downto 0 );
    out_1 : out std_logic_vector( 16-1 downto 0 );
    out_2 : out std_logic_vector( 16-1 downto 0 );
    out_3 : out std_logic_vector( 16-1 downto 0 );
    out_4 : out std_logic_vector( 16-1 downto 0 );
    out_5 : out std_logic_vector( 16-1 downto 0 );
    out_6 : out std_logic_vector( 16-1 downto 0 );
    out_7 : out std_logic_vector( 16-1 downto 0 );
    out_8 : out std_logic_vector( 16-1 downto 0 );
    out_9 : out std_logic_vector( 16-1 downto 0 );
    out_10 : out std_logic_vector( 16-1 downto 0 );
    out_11 : out std_logic_vector( 16-1 downto 0 );
    out_12 : out std_logic_vector( 16-1 downto 0 );
    out_13 : out std_logic_vector( 16-1 downto 0 );
    out_14 : out std_logic_vector( 16-1 downto 0 );
    out_15 : out std_logic_vector( 16-1 downto 0 );
    out_16 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_vector_reinterpret6;
architecture structural of psb3_0_vector_reinterpret6 is 
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 16-1 downto 0 );
begin
  out_1 <= reinterpret0_output_port_net;
  out_2 <= reinterpret1_output_port_net;
  out_3 <= reinterpret2_output_port_net;
  out_4 <= reinterpret3_output_port_net;
  out_5 <= reinterpret4_output_port_net;
  out_6 <= reinterpret5_output_port_net;
  out_7 <= reinterpret6_output_port_net;
  out_8 <= reinterpret7_output_port_net;
  out_9 <= reinterpret8_output_port_net;
  out_10 <= reinterpret9_output_port_net;
  out_11 <= reinterpret10_output_port_net;
  out_12 <= reinterpret11_output_port_net;
  out_13 <= reinterpret12_output_port_net;
  out_14 <= reinterpret13_output_port_net;
  out_15 <= reinterpret14_output_port_net;
  out_16 <= reinterpret15_output_port_net;
  slice0_y_net <= in_1;
  slice1_y_net <= in_2;
  slice2_y_net <= in_3;
  slice3_y_net <= in_4;
  slice4_y_net <= in_5;
  slice5_y_net <= in_6;
  slice6_y_net <= in_7;
  slice7_y_net <= in_8;
  slice8_y_net <= in_9;
  slice9_y_net <= in_10;
  slice10_y_net <= in_11;
  slice11_y_net <= in_12;
  slice12_y_net <= in_13;
  slice13_y_net <= in_14;
  slice14_y_net <= in_15;
  slice15_y_net <= in_16;
  reinterpret0 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice0_y_net,
    output_port => reinterpret0_output_port_net
  );
  reinterpret1 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice1_y_net,
    output_port => reinterpret1_output_port_net
  );
  reinterpret2 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice2_y_net,
    output_port => reinterpret2_output_port_net
  );
  reinterpret3 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice3_y_net,
    output_port => reinterpret3_output_port_net
  );
  reinterpret4 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice4_y_net,
    output_port => reinterpret4_output_port_net
  );
  reinterpret5 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice5_y_net,
    output_port => reinterpret5_output_port_net
  );
  reinterpret6 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice6_y_net,
    output_port => reinterpret6_output_port_net
  );
  reinterpret7 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice7_y_net,
    output_port => reinterpret7_output_port_net
  );
  reinterpret8 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice8_y_net,
    output_port => reinterpret8_output_port_net
  );
  reinterpret9 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice9_y_net,
    output_port => reinterpret9_output_port_net
  );
  reinterpret10 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice10_y_net,
    output_port => reinterpret10_output_port_net
  );
  reinterpret11 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice11_y_net,
    output_port => reinterpret11_output_port_net
  );
  reinterpret12 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice12_y_net,
    output_port => reinterpret12_output_port_net
  );
  reinterpret13 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice13_y_net,
    output_port => reinterpret13_output_port_net
  );
  reinterpret14 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice14_y_net,
    output_port => reinterpret14_output_port_net
  );
  reinterpret15 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice15_y_net,
    output_port => reinterpret15_output_port_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Vector Reinterpret7
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_reinterpret7 is
  port (
    in_1 : in std_logic_vector( 16-1 downto 0 );
    in_2 : in std_logic_vector( 16-1 downto 0 );
    in_3 : in std_logic_vector( 16-1 downto 0 );
    in_4 : in std_logic_vector( 16-1 downto 0 );
    in_5 : in std_logic_vector( 16-1 downto 0 );
    in_6 : in std_logic_vector( 16-1 downto 0 );
    in_7 : in std_logic_vector( 16-1 downto 0 );
    in_8 : in std_logic_vector( 16-1 downto 0 );
    in_9 : in std_logic_vector( 16-1 downto 0 );
    in_10 : in std_logic_vector( 16-1 downto 0 );
    in_11 : in std_logic_vector( 16-1 downto 0 );
    in_12 : in std_logic_vector( 16-1 downto 0 );
    in_13 : in std_logic_vector( 16-1 downto 0 );
    in_14 : in std_logic_vector( 16-1 downto 0 );
    in_15 : in std_logic_vector( 16-1 downto 0 );
    in_16 : in std_logic_vector( 16-1 downto 0 );
    out_1 : out std_logic_vector( 16-1 downto 0 );
    out_2 : out std_logic_vector( 16-1 downto 0 );
    out_3 : out std_logic_vector( 16-1 downto 0 );
    out_4 : out std_logic_vector( 16-1 downto 0 );
    out_5 : out std_logic_vector( 16-1 downto 0 );
    out_6 : out std_logic_vector( 16-1 downto 0 );
    out_7 : out std_logic_vector( 16-1 downto 0 );
    out_8 : out std_logic_vector( 16-1 downto 0 );
    out_9 : out std_logic_vector( 16-1 downto 0 );
    out_10 : out std_logic_vector( 16-1 downto 0 );
    out_11 : out std_logic_vector( 16-1 downto 0 );
    out_12 : out std_logic_vector( 16-1 downto 0 );
    out_13 : out std_logic_vector( 16-1 downto 0 );
    out_14 : out std_logic_vector( 16-1 downto 0 );
    out_15 : out std_logic_vector( 16-1 downto 0 );
    out_16 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_vector_reinterpret7;
architecture structural of psb3_0_vector_reinterpret7 is 
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub8_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub6_s_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub0_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub5_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub10_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub11_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub12_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub13_s_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub14_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub7_s_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub15_s_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub9_s_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub3_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
begin
  out_1 <= reinterpret0_output_port_net;
  out_2 <= reinterpret1_output_port_net;
  out_3 <= reinterpret2_output_port_net;
  out_4 <= reinterpret3_output_port_net;
  out_5 <= reinterpret4_output_port_net;
  out_6 <= reinterpret5_output_port_net;
  out_7 <= reinterpret6_output_port_net;
  out_8 <= reinterpret7_output_port_net;
  out_9 <= reinterpret8_output_port_net;
  out_10 <= reinterpret9_output_port_net;
  out_11 <= reinterpret10_output_port_net;
  out_12 <= reinterpret11_output_port_net;
  out_13 <= reinterpret12_output_port_net;
  out_14 <= reinterpret13_output_port_net;
  out_15 <= reinterpret14_output_port_net;
  out_16 <= reinterpret15_output_port_net;
  addsub0_s_net <= in_1;
  addsub1_s_net <= in_2;
  addsub2_s_net <= in_3;
  addsub3_s_net <= in_4;
  addsub4_s_net <= in_5;
  addsub5_s_net <= in_6;
  addsub6_s_net <= in_7;
  addsub7_s_net <= in_8;
  addsub8_s_net <= in_9;
  addsub9_s_net <= in_10;
  addsub10_s_net <= in_11;
  addsub11_s_net <= in_12;
  addsub12_s_net <= in_13;
  addsub13_s_net <= in_14;
  addsub14_s_net <= in_15;
  addsub15_s_net <= in_16;
  reinterpret0 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub0_s_net,
    output_port => reinterpret0_output_port_net
  );
  reinterpret1 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub1_s_net,
    output_port => reinterpret1_output_port_net
  );
  reinterpret2 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub2_s_net,
    output_port => reinterpret2_output_port_net
  );
  reinterpret3 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub3_s_net,
    output_port => reinterpret3_output_port_net
  );
  reinterpret4 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub4_s_net,
    output_port => reinterpret4_output_port_net
  );
  reinterpret5 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub5_s_net,
    output_port => reinterpret5_output_port_net
  );
  reinterpret6 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub6_s_net,
    output_port => reinterpret6_output_port_net
  );
  reinterpret7 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub7_s_net,
    output_port => reinterpret7_output_port_net
  );
  reinterpret8 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub8_s_net,
    output_port => reinterpret8_output_port_net
  );
  reinterpret9 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub9_s_net,
    output_port => reinterpret9_output_port_net
  );
  reinterpret10 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub10_s_net,
    output_port => reinterpret10_output_port_net
  );
  reinterpret11 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub11_s_net,
    output_port => reinterpret11_output_port_net
  );
  reinterpret12 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub12_s_net,
    output_port => reinterpret12_output_port_net
  );
  reinterpret13 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub13_s_net,
    output_port => reinterpret13_output_port_net
  );
  reinterpret14 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub14_s_net,
    output_port => reinterpret14_output_port_net
  );
  reinterpret15 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub15_s_net,
    output_port => reinterpret15_output_port_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Vector Reinterpret8
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_reinterpret8 is
  port (
    in_1 : in std_logic_vector( 16-1 downto 0 );
    in_2 : in std_logic_vector( 16-1 downto 0 );
    in_3 : in std_logic_vector( 16-1 downto 0 );
    in_4 : in std_logic_vector( 16-1 downto 0 );
    in_5 : in std_logic_vector( 16-1 downto 0 );
    in_6 : in std_logic_vector( 16-1 downto 0 );
    in_7 : in std_logic_vector( 16-1 downto 0 );
    in_8 : in std_logic_vector( 16-1 downto 0 );
    in_9 : in std_logic_vector( 16-1 downto 0 );
    in_10 : in std_logic_vector( 16-1 downto 0 );
    in_11 : in std_logic_vector( 16-1 downto 0 );
    in_12 : in std_logic_vector( 16-1 downto 0 );
    in_13 : in std_logic_vector( 16-1 downto 0 );
    in_14 : in std_logic_vector( 16-1 downto 0 );
    in_15 : in std_logic_vector( 16-1 downto 0 );
    in_16 : in std_logic_vector( 16-1 downto 0 );
    out_1 : out std_logic_vector( 16-1 downto 0 );
    out_2 : out std_logic_vector( 16-1 downto 0 );
    out_3 : out std_logic_vector( 16-1 downto 0 );
    out_4 : out std_logic_vector( 16-1 downto 0 );
    out_5 : out std_logic_vector( 16-1 downto 0 );
    out_6 : out std_logic_vector( 16-1 downto 0 );
    out_7 : out std_logic_vector( 16-1 downto 0 );
    out_8 : out std_logic_vector( 16-1 downto 0 );
    out_9 : out std_logic_vector( 16-1 downto 0 );
    out_10 : out std_logic_vector( 16-1 downto 0 );
    out_11 : out std_logic_vector( 16-1 downto 0 );
    out_12 : out std_logic_vector( 16-1 downto 0 );
    out_13 : out std_logic_vector( 16-1 downto 0 );
    out_14 : out std_logic_vector( 16-1 downto 0 );
    out_15 : out std_logic_vector( 16-1 downto 0 );
    out_16 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_vector_reinterpret8;
architecture structural of psb3_0_vector_reinterpret8 is 
  signal addsub10_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub11_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub12_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub15_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub13_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub14_s_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub7_s_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub8_s_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub9_s_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub0_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal addsub3_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub5_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub6_s_net : std_logic_vector( 16-1 downto 0 );
begin
  out_1 <= reinterpret0_output_port_net;
  out_2 <= reinterpret1_output_port_net;
  out_3 <= reinterpret2_output_port_net;
  out_4 <= reinterpret3_output_port_net;
  out_5 <= reinterpret4_output_port_net;
  out_6 <= reinterpret5_output_port_net;
  out_7 <= reinterpret6_output_port_net;
  out_8 <= reinterpret7_output_port_net;
  out_9 <= reinterpret8_output_port_net;
  out_10 <= reinterpret9_output_port_net;
  out_11 <= reinterpret10_output_port_net;
  out_12 <= reinterpret11_output_port_net;
  out_13 <= reinterpret12_output_port_net;
  out_14 <= reinterpret13_output_port_net;
  out_15 <= reinterpret14_output_port_net;
  out_16 <= reinterpret15_output_port_net;
  addsub0_s_net <= in_1;
  addsub1_s_net <= in_2;
  addsub2_s_net <= in_3;
  addsub3_s_net <= in_4;
  addsub4_s_net <= in_5;
  addsub5_s_net <= in_6;
  addsub6_s_net <= in_7;
  addsub7_s_net <= in_8;
  addsub8_s_net <= in_9;
  addsub9_s_net <= in_10;
  addsub10_s_net <= in_11;
  addsub11_s_net <= in_12;
  addsub12_s_net <= in_13;
  addsub13_s_net <= in_14;
  addsub14_s_net <= in_15;
  addsub15_s_net <= in_16;
  reinterpret0 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub0_s_net,
    output_port => reinterpret0_output_port_net
  );
  reinterpret1 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub1_s_net,
    output_port => reinterpret1_output_port_net
  );
  reinterpret2 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub2_s_net,
    output_port => reinterpret2_output_port_net
  );
  reinterpret3 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub3_s_net,
    output_port => reinterpret3_output_port_net
  );
  reinterpret4 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub4_s_net,
    output_port => reinterpret4_output_port_net
  );
  reinterpret5 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub5_s_net,
    output_port => reinterpret5_output_port_net
  );
  reinterpret6 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub6_s_net,
    output_port => reinterpret6_output_port_net
  );
  reinterpret7 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub7_s_net,
    output_port => reinterpret7_output_port_net
  );
  reinterpret8 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub8_s_net,
    output_port => reinterpret8_output_port_net
  );
  reinterpret9 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub9_s_net,
    output_port => reinterpret9_output_port_net
  );
  reinterpret10 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub10_s_net,
    output_port => reinterpret10_output_port_net
  );
  reinterpret11 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub11_s_net,
    output_port => reinterpret11_output_port_net
  );
  reinterpret12 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub12_s_net,
    output_port => reinterpret12_output_port_net
  );
  reinterpret13 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub13_s_net,
    output_port => reinterpret13_output_port_net
  );
  reinterpret14 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub14_s_net,
    output_port => reinterpret14_output_port_net
  );
  reinterpret15 : entity xil_defaultlib.sysgen_reinterpret_2d4abf6691 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => addsub15_s_net,
    output_port => reinterpret15_output_port_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Vector Reinterpret9
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_reinterpret9 is
  port (
    in_1 : in std_logic_vector( 16-1 downto 0 );
    in_2 : in std_logic_vector( 16-1 downto 0 );
    in_3 : in std_logic_vector( 16-1 downto 0 );
    in_4 : in std_logic_vector( 16-1 downto 0 );
    in_5 : in std_logic_vector( 16-1 downto 0 );
    in_6 : in std_logic_vector( 16-1 downto 0 );
    in_7 : in std_logic_vector( 16-1 downto 0 );
    in_8 : in std_logic_vector( 16-1 downto 0 );
    in_9 : in std_logic_vector( 16-1 downto 0 );
    in_10 : in std_logic_vector( 16-1 downto 0 );
    in_11 : in std_logic_vector( 16-1 downto 0 );
    in_12 : in std_logic_vector( 16-1 downto 0 );
    in_13 : in std_logic_vector( 16-1 downto 0 );
    in_14 : in std_logic_vector( 16-1 downto 0 );
    in_15 : in std_logic_vector( 16-1 downto 0 );
    in_16 : in std_logic_vector( 16-1 downto 0 );
    out_1 : out std_logic_vector( 16-1 downto 0 );
    out_2 : out std_logic_vector( 16-1 downto 0 );
    out_3 : out std_logic_vector( 16-1 downto 0 );
    out_4 : out std_logic_vector( 16-1 downto 0 );
    out_5 : out std_logic_vector( 16-1 downto 0 );
    out_6 : out std_logic_vector( 16-1 downto 0 );
    out_7 : out std_logic_vector( 16-1 downto 0 );
    out_8 : out std_logic_vector( 16-1 downto 0 );
    out_9 : out std_logic_vector( 16-1 downto 0 );
    out_10 : out std_logic_vector( 16-1 downto 0 );
    out_11 : out std_logic_vector( 16-1 downto 0 );
    out_12 : out std_logic_vector( 16-1 downto 0 );
    out_13 : out std_logic_vector( 16-1 downto 0 );
    out_14 : out std_logic_vector( 16-1 downto 0 );
    out_15 : out std_logic_vector( 16-1 downto 0 );
    out_16 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_vector_reinterpret9;
architecture structural of psb3_0_vector_reinterpret9 is 
  signal slice1_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 16-1 downto 0 );
begin
  out_1 <= reinterpret0_output_port_net;
  out_2 <= reinterpret1_output_port_net;
  out_3 <= reinterpret2_output_port_net;
  out_4 <= reinterpret3_output_port_net;
  out_5 <= reinterpret4_output_port_net;
  out_6 <= reinterpret5_output_port_net;
  out_7 <= reinterpret6_output_port_net;
  out_8 <= reinterpret7_output_port_net;
  out_9 <= reinterpret8_output_port_net;
  out_10 <= reinterpret9_output_port_net;
  out_11 <= reinterpret10_output_port_net;
  out_12 <= reinterpret11_output_port_net;
  out_13 <= reinterpret12_output_port_net;
  out_14 <= reinterpret13_output_port_net;
  out_15 <= reinterpret14_output_port_net;
  out_16 <= reinterpret15_output_port_net;
  slice0_y_net <= in_1;
  slice1_y_net <= in_2;
  slice2_y_net <= in_3;
  slice3_y_net <= in_4;
  slice4_y_net <= in_5;
  slice5_y_net <= in_6;
  slice6_y_net <= in_7;
  slice7_y_net <= in_8;
  slice8_y_net <= in_9;
  slice9_y_net <= in_10;
  slice10_y_net <= in_11;
  slice11_y_net <= in_12;
  slice12_y_net <= in_13;
  slice13_y_net <= in_14;
  slice14_y_net <= in_15;
  slice15_y_net <= in_16;
  reinterpret0 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice0_y_net,
    output_port => reinterpret0_output_port_net
  );
  reinterpret1 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice1_y_net,
    output_port => reinterpret1_output_port_net
  );
  reinterpret2 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice2_y_net,
    output_port => reinterpret2_output_port_net
  );
  reinterpret3 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice3_y_net,
    output_port => reinterpret3_output_port_net
  );
  reinterpret4 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice4_y_net,
    output_port => reinterpret4_output_port_net
  );
  reinterpret5 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice5_y_net,
    output_port => reinterpret5_output_port_net
  );
  reinterpret6 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice6_y_net,
    output_port => reinterpret6_output_port_net
  );
  reinterpret7 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice7_y_net,
    output_port => reinterpret7_output_port_net
  );
  reinterpret8 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice8_y_net,
    output_port => reinterpret8_output_port_net
  );
  reinterpret9 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice9_y_net,
    output_port => reinterpret9_output_port_net
  );
  reinterpret10 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice10_y_net,
    output_port => reinterpret10_output_port_net
  );
  reinterpret11 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice11_y_net,
    output_port => reinterpret11_output_port_net
  );
  reinterpret12 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice12_y_net,
    output_port => reinterpret12_output_port_net
  );
  reinterpret13 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice13_y_net,
    output_port => reinterpret13_output_port_net
  );
  reinterpret14 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice14_y_net,
    output_port => reinterpret14_output_port_net
  );
  reinterpret15 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice15_y_net,
    output_port => reinterpret15_output_port_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Vector to Scalar
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_to_scalar_x7 is
  port (
    i_1 : in std_logic_vector( 16-1 downto 0 );
    i_2 : in std_logic_vector( 16-1 downto 0 );
    i_3 : in std_logic_vector( 16-1 downto 0 );
    i_4 : in std_logic_vector( 16-1 downto 0 );
    i_5 : in std_logic_vector( 16-1 downto 0 );
    i_6 : in std_logic_vector( 16-1 downto 0 );
    i_7 : in std_logic_vector( 16-1 downto 0 );
    i_8 : in std_logic_vector( 16-1 downto 0 );
    i_9 : in std_logic_vector( 16-1 downto 0 );
    i_10 : in std_logic_vector( 16-1 downto 0 );
    i_11 : in std_logic_vector( 16-1 downto 0 );
    i_12 : in std_logic_vector( 16-1 downto 0 );
    i_13 : in std_logic_vector( 16-1 downto 0 );
    i_14 : in std_logic_vector( 16-1 downto 0 );
    i_15 : in std_logic_vector( 16-1 downto 0 );
    i_16 : in std_logic_vector( 16-1 downto 0 );
    o : out std_logic_vector( 256-1 downto 0 )
  );
end psb3_0_vector_to_scalar_x7;
architecture structural of psb3_0_vector_to_scalar_x7 is 
  signal concat1_y_net : std_logic_vector( 256-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
begin
  o <= concat1_y_net;
  reinterpret0_output_port_net <= i_1;
  reinterpret1_output_port_net <= i_2;
  reinterpret2_output_port_net <= i_3;
  reinterpret3_output_port_net <= i_4;
  reinterpret4_output_port_net <= i_5;
  reinterpret5_output_port_net <= i_6;
  reinterpret6_output_port_net <= i_7;
  reinterpret7_output_port_net <= i_8;
  reinterpret8_output_port_net <= i_9;
  reinterpret9_output_port_net <= i_10;
  reinterpret10_output_port_net <= i_11;
  reinterpret11_output_port_net <= i_12;
  reinterpret12_output_port_net <= i_13;
  reinterpret13_output_port_net <= i_14;
  reinterpret14_output_port_net <= i_15;
  reinterpret15_output_port_net <= i_16;
  concat1 : entity xil_defaultlib.sysgen_concat_6c8db818fa 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => reinterpret15_output_port_net,
    in1 => reinterpret14_output_port_net,
    in2 => reinterpret13_output_port_net,
    in3 => reinterpret12_output_port_net,
    in4 => reinterpret11_output_port_net,
    in5 => reinterpret10_output_port_net,
    in6 => reinterpret9_output_port_net,
    in7 => reinterpret8_output_port_net,
    in8 => reinterpret7_output_port_net,
    in9 => reinterpret6_output_port_net,
    in10 => reinterpret5_output_port_net,
    in11 => reinterpret4_output_port_net,
    in12 => reinterpret3_output_port_net,
    in13 => reinterpret2_output_port_net,
    in14 => reinterpret1_output_port_net,
    in15 => reinterpret0_output_port_net,
    y => concat1_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Vector to Scalar1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_to_scalar1_x7 is
  port (
    i_1 : in std_logic_vector( 16-1 downto 0 );
    i_2 : in std_logic_vector( 16-1 downto 0 );
    i_3 : in std_logic_vector( 16-1 downto 0 );
    i_4 : in std_logic_vector( 16-1 downto 0 );
    i_5 : in std_logic_vector( 16-1 downto 0 );
    i_6 : in std_logic_vector( 16-1 downto 0 );
    i_7 : in std_logic_vector( 16-1 downto 0 );
    i_8 : in std_logic_vector( 16-1 downto 0 );
    i_9 : in std_logic_vector( 16-1 downto 0 );
    i_10 : in std_logic_vector( 16-1 downto 0 );
    i_11 : in std_logic_vector( 16-1 downto 0 );
    i_12 : in std_logic_vector( 16-1 downto 0 );
    i_13 : in std_logic_vector( 16-1 downto 0 );
    i_14 : in std_logic_vector( 16-1 downto 0 );
    i_15 : in std_logic_vector( 16-1 downto 0 );
    i_16 : in std_logic_vector( 16-1 downto 0 );
    o : out std_logic_vector( 256-1 downto 0 )
  );
end psb3_0_vector_to_scalar1_x7;
architecture structural of psb3_0_vector_to_scalar1_x7 is 
  signal concat1_y_net : std_logic_vector( 256-1 downto 0 );
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
begin
  o <= concat1_y_net;
  reinterpret0_output_port_net <= i_1;
  reinterpret1_output_port_net <= i_2;
  reinterpret2_output_port_net <= i_3;
  reinterpret3_output_port_net <= i_4;
  reinterpret4_output_port_net <= i_5;
  reinterpret5_output_port_net <= i_6;
  reinterpret6_output_port_net <= i_7;
  reinterpret7_output_port_net <= i_8;
  reinterpret8_output_port_net <= i_9;
  reinterpret9_output_port_net <= i_10;
  reinterpret10_output_port_net <= i_11;
  reinterpret11_output_port_net <= i_12;
  reinterpret12_output_port_net <= i_13;
  reinterpret13_output_port_net <= i_14;
  reinterpret14_output_port_net <= i_15;
  reinterpret15_output_port_net <= i_16;
  concat1 : entity xil_defaultlib.sysgen_concat_6c8db818fa 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => reinterpret15_output_port_net,
    in1 => reinterpret14_output_port_net,
    in2 => reinterpret13_output_port_net,
    in3 => reinterpret12_output_port_net,
    in4 => reinterpret11_output_port_net,
    in5 => reinterpret10_output_port_net,
    in6 => reinterpret9_output_port_net,
    in7 => reinterpret8_output_port_net,
    in8 => reinterpret7_output_port_net,
    in9 => reinterpret6_output_port_net,
    in10 => reinterpret5_output_port_net,
    in11 => reinterpret4_output_port_net,
    in12 => reinterpret3_output_port_net,
    in13 => reinterpret2_output_port_net,
    in14 => reinterpret1_output_port_net,
    in15 => reinterpret0_output_port_net,
    y => concat1_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Vector to Scalar2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_to_scalar2_x7 is
  port (
    i_1 : in std_logic_vector( 16-1 downto 0 );
    i_2 : in std_logic_vector( 16-1 downto 0 );
    i_3 : in std_logic_vector( 16-1 downto 0 );
    i_4 : in std_logic_vector( 16-1 downto 0 );
    i_5 : in std_logic_vector( 16-1 downto 0 );
    i_6 : in std_logic_vector( 16-1 downto 0 );
    i_7 : in std_logic_vector( 16-1 downto 0 );
    i_8 : in std_logic_vector( 16-1 downto 0 );
    i_9 : in std_logic_vector( 16-1 downto 0 );
    i_10 : in std_logic_vector( 16-1 downto 0 );
    i_11 : in std_logic_vector( 16-1 downto 0 );
    i_12 : in std_logic_vector( 16-1 downto 0 );
    i_13 : in std_logic_vector( 16-1 downto 0 );
    i_14 : in std_logic_vector( 16-1 downto 0 );
    i_15 : in std_logic_vector( 16-1 downto 0 );
    i_16 : in std_logic_vector( 16-1 downto 0 );
    o : out std_logic_vector( 256-1 downto 0 )
  );
end psb3_0_vector_to_scalar2_x7;
architecture structural of psb3_0_vector_to_scalar2_x7 is 
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal concat1_y_net : std_logic_vector( 256-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
begin
  o <= concat1_y_net;
  reinterpret0_output_port_net <= i_1;
  reinterpret1_output_port_net <= i_2;
  reinterpret2_output_port_net <= i_3;
  reinterpret3_output_port_net <= i_4;
  reinterpret4_output_port_net <= i_5;
  reinterpret5_output_port_net <= i_6;
  reinterpret6_output_port_net <= i_7;
  reinterpret7_output_port_net <= i_8;
  reinterpret8_output_port_net <= i_9;
  reinterpret9_output_port_net <= i_10;
  reinterpret10_output_port_net <= i_11;
  reinterpret11_output_port_net <= i_12;
  reinterpret12_output_port_net <= i_13;
  reinterpret13_output_port_net <= i_14;
  reinterpret14_output_port_net <= i_15;
  reinterpret15_output_port_net <= i_16;
  concat1 : entity xil_defaultlib.sysgen_concat_6c8db818fa 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => reinterpret15_output_port_net,
    in1 => reinterpret14_output_port_net,
    in2 => reinterpret13_output_port_net,
    in3 => reinterpret12_output_port_net,
    in4 => reinterpret11_output_port_net,
    in5 => reinterpret10_output_port_net,
    in6 => reinterpret9_output_port_net,
    in7 => reinterpret8_output_port_net,
    in8 => reinterpret7_output_port_net,
    in9 => reinterpret6_output_port_net,
    in10 => reinterpret5_output_port_net,
    in11 => reinterpret4_output_port_net,
    in12 => reinterpret3_output_port_net,
    in13 => reinterpret2_output_port_net,
    in14 => reinterpret1_output_port_net,
    in15 => reinterpret0_output_port_net,
    y => concat1_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Vector to Scalar3
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_to_scalar3 is
  port (
    i_1 : in std_logic_vector( 16-1 downto 0 );
    i_2 : in std_logic_vector( 16-1 downto 0 );
    i_3 : in std_logic_vector( 16-1 downto 0 );
    i_4 : in std_logic_vector( 16-1 downto 0 );
    i_5 : in std_logic_vector( 16-1 downto 0 );
    i_6 : in std_logic_vector( 16-1 downto 0 );
    i_7 : in std_logic_vector( 16-1 downto 0 );
    i_8 : in std_logic_vector( 16-1 downto 0 );
    i_9 : in std_logic_vector( 16-1 downto 0 );
    i_10 : in std_logic_vector( 16-1 downto 0 );
    i_11 : in std_logic_vector( 16-1 downto 0 );
    i_12 : in std_logic_vector( 16-1 downto 0 );
    i_13 : in std_logic_vector( 16-1 downto 0 );
    i_14 : in std_logic_vector( 16-1 downto 0 );
    i_15 : in std_logic_vector( 16-1 downto 0 );
    i_16 : in std_logic_vector( 16-1 downto 0 );
    o : out std_logic_vector( 256-1 downto 0 )
  );
end psb3_0_vector_to_scalar3;
architecture structural of psb3_0_vector_to_scalar3 is 
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal concat1_y_net : std_logic_vector( 256-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
begin
  o <= concat1_y_net;
  reinterpret0_output_port_net <= i_1;
  reinterpret1_output_port_net <= i_2;
  reinterpret2_output_port_net <= i_3;
  reinterpret3_output_port_net <= i_4;
  reinterpret4_output_port_net <= i_5;
  reinterpret5_output_port_net <= i_6;
  reinterpret6_output_port_net <= i_7;
  reinterpret7_output_port_net <= i_8;
  reinterpret8_output_port_net <= i_9;
  reinterpret9_output_port_net <= i_10;
  reinterpret10_output_port_net <= i_11;
  reinterpret11_output_port_net <= i_12;
  reinterpret12_output_port_net <= i_13;
  reinterpret13_output_port_net <= i_14;
  reinterpret14_output_port_net <= i_15;
  reinterpret15_output_port_net <= i_16;
  concat1 : entity xil_defaultlib.sysgen_concat_6c8db818fa 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => reinterpret15_output_port_net,
    in1 => reinterpret14_output_port_net,
    in2 => reinterpret13_output_port_net,
    in3 => reinterpret12_output_port_net,
    in4 => reinterpret11_output_port_net,
    in5 => reinterpret10_output_port_net,
    in6 => reinterpret9_output_port_net,
    in7 => reinterpret8_output_port_net,
    in8 => reinterpret7_output_port_net,
    in9 => reinterpret6_output_port_net,
    in10 => reinterpret5_output_port_net,
    in11 => reinterpret4_output_port_net,
    in12 => reinterpret3_output_port_net,
    in13 => reinterpret2_output_port_net,
    in14 => reinterpret1_output_port_net,
    in15 => reinterpret0_output_port_net,
    y => concat1_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Vector to Scalar4
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_to_scalar4 is
  port (
    i_1 : in std_logic_vector( 16-1 downto 0 );
    i_2 : in std_logic_vector( 16-1 downto 0 );
    i_3 : in std_logic_vector( 16-1 downto 0 );
    i_4 : in std_logic_vector( 16-1 downto 0 );
    i_5 : in std_logic_vector( 16-1 downto 0 );
    i_6 : in std_logic_vector( 16-1 downto 0 );
    i_7 : in std_logic_vector( 16-1 downto 0 );
    i_8 : in std_logic_vector( 16-1 downto 0 );
    i_9 : in std_logic_vector( 16-1 downto 0 );
    i_10 : in std_logic_vector( 16-1 downto 0 );
    i_11 : in std_logic_vector( 16-1 downto 0 );
    i_12 : in std_logic_vector( 16-1 downto 0 );
    i_13 : in std_logic_vector( 16-1 downto 0 );
    i_14 : in std_logic_vector( 16-1 downto 0 );
    i_15 : in std_logic_vector( 16-1 downto 0 );
    i_16 : in std_logic_vector( 16-1 downto 0 );
    o : out std_logic_vector( 256-1 downto 0 )
  );
end psb3_0_vector_to_scalar4;
architecture structural of psb3_0_vector_to_scalar4 is 
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal concat1_y_net : std_logic_vector( 256-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
begin
  o <= concat1_y_net;
  reinterpret0_output_port_net <= i_1;
  reinterpret1_output_port_net <= i_2;
  reinterpret2_output_port_net <= i_3;
  reinterpret3_output_port_net <= i_4;
  reinterpret4_output_port_net <= i_5;
  reinterpret5_output_port_net <= i_6;
  reinterpret6_output_port_net <= i_7;
  reinterpret7_output_port_net <= i_8;
  reinterpret8_output_port_net <= i_9;
  reinterpret9_output_port_net <= i_10;
  reinterpret10_output_port_net <= i_11;
  reinterpret11_output_port_net <= i_12;
  reinterpret12_output_port_net <= i_13;
  reinterpret13_output_port_net <= i_14;
  reinterpret14_output_port_net <= i_15;
  reinterpret15_output_port_net <= i_16;
  concat1 : entity xil_defaultlib.sysgen_concat_6c8db818fa 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => reinterpret15_output_port_net,
    in1 => reinterpret14_output_port_net,
    in2 => reinterpret13_output_port_net,
    in3 => reinterpret12_output_port_net,
    in4 => reinterpret11_output_port_net,
    in5 => reinterpret10_output_port_net,
    in6 => reinterpret9_output_port_net,
    in7 => reinterpret8_output_port_net,
    in8 => reinterpret7_output_port_net,
    in9 => reinterpret6_output_port_net,
    in10 => reinterpret5_output_port_net,
    in11 => reinterpret4_output_port_net,
    in12 => reinterpret3_output_port_net,
    in13 => reinterpret2_output_port_net,
    in14 => reinterpret1_output_port_net,
    in15 => reinterpret0_output_port_net,
    y => concat1_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Vector to Scalar5
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_to_scalar5 is
  port (
    i_1 : in std_logic_vector( 16-1 downto 0 );
    i_2 : in std_logic_vector( 16-1 downto 0 );
    i_3 : in std_logic_vector( 16-1 downto 0 );
    i_4 : in std_logic_vector( 16-1 downto 0 );
    i_5 : in std_logic_vector( 16-1 downto 0 );
    i_6 : in std_logic_vector( 16-1 downto 0 );
    i_7 : in std_logic_vector( 16-1 downto 0 );
    i_8 : in std_logic_vector( 16-1 downto 0 );
    i_9 : in std_logic_vector( 16-1 downto 0 );
    i_10 : in std_logic_vector( 16-1 downto 0 );
    i_11 : in std_logic_vector( 16-1 downto 0 );
    i_12 : in std_logic_vector( 16-1 downto 0 );
    i_13 : in std_logic_vector( 16-1 downto 0 );
    i_14 : in std_logic_vector( 16-1 downto 0 );
    i_15 : in std_logic_vector( 16-1 downto 0 );
    i_16 : in std_logic_vector( 16-1 downto 0 );
    o : out std_logic_vector( 256-1 downto 0 )
  );
end psb3_0_vector_to_scalar5;
architecture structural of psb3_0_vector_to_scalar5 is 
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal concat1_y_net : std_logic_vector( 256-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
begin
  o <= concat1_y_net;
  reinterpret0_output_port_net <= i_1;
  reinterpret1_output_port_net <= i_2;
  reinterpret2_output_port_net <= i_3;
  reinterpret3_output_port_net <= i_4;
  reinterpret4_output_port_net <= i_5;
  reinterpret5_output_port_net <= i_6;
  reinterpret6_output_port_net <= i_7;
  reinterpret7_output_port_net <= i_8;
  reinterpret8_output_port_net <= i_9;
  reinterpret9_output_port_net <= i_10;
  reinterpret10_output_port_net <= i_11;
  reinterpret11_output_port_net <= i_12;
  reinterpret12_output_port_net <= i_13;
  reinterpret13_output_port_net <= i_14;
  reinterpret14_output_port_net <= i_15;
  reinterpret15_output_port_net <= i_16;
  concat1 : entity xil_defaultlib.sysgen_concat_6c8db818fa 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => reinterpret15_output_port_net,
    in1 => reinterpret14_output_port_net,
    in2 => reinterpret13_output_port_net,
    in3 => reinterpret12_output_port_net,
    in4 => reinterpret11_output_port_net,
    in5 => reinterpret10_output_port_net,
    in6 => reinterpret9_output_port_net,
    in7 => reinterpret8_output_port_net,
    in8 => reinterpret7_output_port_net,
    in9 => reinterpret6_output_port_net,
    in10 => reinterpret5_output_port_net,
    in11 => reinterpret4_output_port_net,
    in12 => reinterpret3_output_port_net,
    in13 => reinterpret2_output_port_net,
    in14 => reinterpret1_output_port_net,
    in15 => reinterpret0_output_port_net,
    y => concat1_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Vector to Scalar6
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_to_scalar6 is
  port (
    i_1 : in std_logic_vector( 16-1 downto 0 );
    i_2 : in std_logic_vector( 16-1 downto 0 );
    i_3 : in std_logic_vector( 16-1 downto 0 );
    i_4 : in std_logic_vector( 16-1 downto 0 );
    i_5 : in std_logic_vector( 16-1 downto 0 );
    i_6 : in std_logic_vector( 16-1 downto 0 );
    i_7 : in std_logic_vector( 16-1 downto 0 );
    i_8 : in std_logic_vector( 16-1 downto 0 );
    i_9 : in std_logic_vector( 16-1 downto 0 );
    i_10 : in std_logic_vector( 16-1 downto 0 );
    i_11 : in std_logic_vector( 16-1 downto 0 );
    i_12 : in std_logic_vector( 16-1 downto 0 );
    i_13 : in std_logic_vector( 16-1 downto 0 );
    i_14 : in std_logic_vector( 16-1 downto 0 );
    i_15 : in std_logic_vector( 16-1 downto 0 );
    i_16 : in std_logic_vector( 16-1 downto 0 );
    o : out std_logic_vector( 256-1 downto 0 )
  );
end psb3_0_vector_to_scalar6;
architecture structural of psb3_0_vector_to_scalar6 is 
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal concat1_y_net : std_logic_vector( 256-1 downto 0 );
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
begin
  o <= concat1_y_net;
  reinterpret0_output_port_net <= i_1;
  reinterpret1_output_port_net <= i_2;
  reinterpret2_output_port_net <= i_3;
  reinterpret3_output_port_net <= i_4;
  reinterpret4_output_port_net <= i_5;
  reinterpret5_output_port_net <= i_6;
  reinterpret6_output_port_net <= i_7;
  reinterpret7_output_port_net <= i_8;
  reinterpret8_output_port_net <= i_9;
  reinterpret9_output_port_net <= i_10;
  reinterpret10_output_port_net <= i_11;
  reinterpret11_output_port_net <= i_12;
  reinterpret12_output_port_net <= i_13;
  reinterpret13_output_port_net <= i_14;
  reinterpret14_output_port_net <= i_15;
  reinterpret15_output_port_net <= i_16;
  concat1 : entity xil_defaultlib.sysgen_concat_6c8db818fa 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => reinterpret15_output_port_net,
    in1 => reinterpret14_output_port_net,
    in2 => reinterpret13_output_port_net,
    in3 => reinterpret12_output_port_net,
    in4 => reinterpret11_output_port_net,
    in5 => reinterpret10_output_port_net,
    in6 => reinterpret9_output_port_net,
    in7 => reinterpret8_output_port_net,
    in8 => reinterpret7_output_port_net,
    in9 => reinterpret6_output_port_net,
    in10 => reinterpret5_output_port_net,
    in11 => reinterpret4_output_port_net,
    in12 => reinterpret3_output_port_net,
    in13 => reinterpret2_output_port_net,
    in14 => reinterpret1_output_port_net,
    in15 => reinterpret0_output_port_net,
    y => concat1_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/Vector to Scalar7
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_to_scalar7 is
  port (
    i_1 : in std_logic_vector( 16-1 downto 0 );
    i_2 : in std_logic_vector( 16-1 downto 0 );
    i_3 : in std_logic_vector( 16-1 downto 0 );
    i_4 : in std_logic_vector( 16-1 downto 0 );
    i_5 : in std_logic_vector( 16-1 downto 0 );
    i_6 : in std_logic_vector( 16-1 downto 0 );
    i_7 : in std_logic_vector( 16-1 downto 0 );
    i_8 : in std_logic_vector( 16-1 downto 0 );
    i_9 : in std_logic_vector( 16-1 downto 0 );
    i_10 : in std_logic_vector( 16-1 downto 0 );
    i_11 : in std_logic_vector( 16-1 downto 0 );
    i_12 : in std_logic_vector( 16-1 downto 0 );
    i_13 : in std_logic_vector( 16-1 downto 0 );
    i_14 : in std_logic_vector( 16-1 downto 0 );
    i_15 : in std_logic_vector( 16-1 downto 0 );
    i_16 : in std_logic_vector( 16-1 downto 0 );
    o : out std_logic_vector( 256-1 downto 0 )
  );
end psb3_0_vector_to_scalar7;
architecture structural of psb3_0_vector_to_scalar7 is 
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal concat1_y_net : std_logic_vector( 256-1 downto 0 );
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
begin
  o <= concat1_y_net;
  reinterpret0_output_port_net <= i_1;
  reinterpret1_output_port_net <= i_2;
  reinterpret2_output_port_net <= i_3;
  reinterpret3_output_port_net <= i_4;
  reinterpret4_output_port_net <= i_5;
  reinterpret5_output_port_net <= i_6;
  reinterpret6_output_port_net <= i_7;
  reinterpret7_output_port_net <= i_8;
  reinterpret8_output_port_net <= i_9;
  reinterpret9_output_port_net <= i_10;
  reinterpret10_output_port_net <= i_11;
  reinterpret11_output_port_net <= i_12;
  reinterpret12_output_port_net <= i_13;
  reinterpret13_output_port_net <= i_14;
  reinterpret14_output_port_net <= i_15;
  reinterpret15_output_port_net <= i_16;
  concat1 : entity xil_defaultlib.sysgen_concat_6c8db818fa 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => reinterpret15_output_port_net,
    in1 => reinterpret14_output_port_net,
    in2 => reinterpret13_output_port_net,
    in3 => reinterpret12_output_port_net,
    in4 => reinterpret11_output_port_net,
    in5 => reinterpret10_output_port_net,
    in6 => reinterpret9_output_port_net,
    in7 => reinterpret8_output_port_net,
    in8 => reinterpret7_output_port_net,
    in9 => reinterpret6_output_port_net,
    in10 => reinterpret5_output_port_net,
    in11 => reinterpret4_output_port_net,
    in12 => reinterpret3_output_port_net,
    in13 => reinterpret2_output_port_net,
    in14 => reinterpret1_output_port_net,
    in15 => reinterpret0_output_port_net,
    y => concat1_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/delayCounter
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_delaycounter is
  port (
    edge1 : in std_logic_vector( 1-1 downto 0 );
    edge2 : in std_logic;
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    delay : out std_logic_vector( 12-1 downto 0 )
  );
end psb3_0_delaycounter;
architecture structural of psb3_0_delaycounter is 
  signal counter1_op_net : std_logic_vector( 12-1 downto 0 );
  signal ce_net : std_logic;
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
  signal register1_q_net : std_logic_vector( 1-1 downto 0 );
  signal register2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay11_q_net : std_logic_vector( 1-1 downto 0 );
  signal test_systolicfft_vhdl_black_box_vo_net : std_logic;
  signal clk_net : std_logic;
  signal const1_op_net : std_logic_vector( 1-1 downto 0 );
begin
  delay <= counter1_op_net;
  delay11_q_net <= edge1;
  test_systolicfft_vhdl_black_box_vo_net <= edge2;
  clk_net <= clk_1;
  ce_net <= ce_1;
  counter1 : entity xil_defaultlib.psb3_0_xlcounter_free 
  generic map (
    core_name0 => "psb3_0_c_counter_binary_v12_0_i2",
    op_arith => xlUnsigned,
    op_width => 12
  )
  port map (
    rst => "0",
    clr => '0',
    en => logical_y_net,
    clk => clk_net,
    ce => ce_net,
    op => counter1_op_net
  );
  logical : entity xil_defaultlib.sysgen_logical_e072b658e1 
  port map (
    clr => '0',
    d0 => register1_q_net,
    d1 => register2_q_net,
    clk => clk_net,
    ce => ce_net,
    y => logical_y_net
  );
  register1 : entity xil_defaultlib.psb3_0_xlregister 
  generic map (
    d_width => 1,
    init_value => b"0"
  )
  port map (
    rst => "0",
    d => const1_op_net,
    en => delay11_q_net,
    clk => clk_net,
    ce => ce_net,
    q => register1_q_net
  );
  register2 : entity xil_defaultlib.psb3_0_xlregister 
  generic map (
    d_width => 1,
    init_value => b"0"
  )
  port map (
    rst => "0",
    d => const1_op_net,
    en(0) => test_systolicfft_vhdl_black_box_vo_net,
    clk => clk_net,
    ce => ce_net,
    q => register2_q_net
  );
  const1 : entity xil_defaultlib.sysgen_constant_71e89d757c 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => const1_op_net
  );
end structural;
-- Generated from Simulink block PSB3_0/ov_detector_IFFT_im/Vector Absolute
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_absolute is
  port (
    d_1 : in std_logic_vector( 20-1 downto 0 );
    d_2 : in std_logic_vector( 20-1 downto 0 );
    d_3 : in std_logic_vector( 20-1 downto 0 );
    d_4 : in std_logic_vector( 20-1 downto 0 );
    d_5 : in std_logic_vector( 20-1 downto 0 );
    d_6 : in std_logic_vector( 20-1 downto 0 );
    d_7 : in std_logic_vector( 20-1 downto 0 );
    d_8 : in std_logic_vector( 20-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    q_1 : out std_logic_vector( 20-1 downto 0 );
    q_2 : out std_logic_vector( 20-1 downto 0 );
    q_3 : out std_logic_vector( 20-1 downto 0 );
    q_4 : out std_logic_vector( 20-1 downto 0 );
    q_5 : out std_logic_vector( 20-1 downto 0 );
    q_6 : out std_logic_vector( 20-1 downto 0 );
    q_7 : out std_logic_vector( 20-1 downto 0 );
    q_8 : out std_logic_vector( 20-1 downto 0 )
  );
end psb3_0_vector_absolute;
architecture structural of psb3_0_vector_absolute is 
  signal ce_net : std_logic;
  signal absolute7_op_net : std_logic_vector( 20-1 downto 0 );
  signal absolute5_op_net : std_logic_vector( 20-1 downto 0 );
  signal clk_net : std_logic;
  signal absolute2_op_net : std_logic_vector( 20-1 downto 0 );
  signal absolute0_op_net : std_logic_vector( 20-1 downto 0 );
  signal absolute6_op_net : std_logic_vector( 20-1 downto 0 );
  signal register0_q_net : std_logic_vector( 20-1 downto 0 );
  signal absolute4_op_net : std_logic_vector( 20-1 downto 0 );
  signal register3_q_net : std_logic_vector( 20-1 downto 0 );
  signal register2_q_net : std_logic_vector( 20-1 downto 0 );
  signal register4_q_net : std_logic_vector( 20-1 downto 0 );
  signal register7_q_net : std_logic_vector( 20-1 downto 0 );
  signal register5_q_net : std_logic_vector( 20-1 downto 0 );
  signal absolute1_op_net : std_logic_vector( 20-1 downto 0 );
  signal absolute3_op_net : std_logic_vector( 20-1 downto 0 );
  signal register1_q_net : std_logic_vector( 20-1 downto 0 );
  signal register6_q_net : std_logic_vector( 20-1 downto 0 );
begin
  q_1 <= absolute0_op_net;
  q_2 <= absolute1_op_net;
  q_3 <= absolute2_op_net;
  q_4 <= absolute3_op_net;
  q_5 <= absolute4_op_net;
  q_6 <= absolute5_op_net;
  q_7 <= absolute6_op_net;
  q_8 <= absolute7_op_net;
  register0_q_net <= d_1;
  register1_q_net <= d_2;
  register2_q_net <= d_3;
  register3_q_net <= d_4;
  register4_q_net <= d_5;
  register5_q_net <= d_6;
  register6_q_net <= d_7;
  register7_q_net <= d_8;
  clk_net <= clk_1;
  ce_net <= ce_1;
  absolute0 : entity xil_defaultlib.sysgen_abs_0161aa1824 
  port map (
    clr => '0',
    a => register0_q_net,
    clk => clk_net,
    ce => ce_net,
    op => absolute0_op_net
  );
  absolute1 : entity xil_defaultlib.sysgen_abs_0161aa1824 
  port map (
    clr => '0',
    a => register1_q_net,
    clk => clk_net,
    ce => ce_net,
    op => absolute1_op_net
  );
  absolute2 : entity xil_defaultlib.sysgen_abs_0161aa1824 
  port map (
    clr => '0',
    a => register2_q_net,
    clk => clk_net,
    ce => ce_net,
    op => absolute2_op_net
  );
  absolute3 : entity xil_defaultlib.sysgen_abs_0161aa1824 
  port map (
    clr => '0',
    a => register3_q_net,
    clk => clk_net,
    ce => ce_net,
    op => absolute3_op_net
  );
  absolute4 : entity xil_defaultlib.sysgen_abs_0161aa1824 
  port map (
    clr => '0',
    a => register4_q_net,
    clk => clk_net,
    ce => ce_net,
    op => absolute4_op_net
  );
  absolute5 : entity xil_defaultlib.sysgen_abs_0161aa1824 
  port map (
    clr => '0',
    a => register5_q_net,
    clk => clk_net,
    ce => ce_net,
    op => absolute5_op_net
  );
  absolute6 : entity xil_defaultlib.sysgen_abs_0161aa1824 
  port map (
    clr => '0',
    a => register6_q_net,
    clk => clk_net,
    ce => ce_net,
    op => absolute6_op_net
  );
  absolute7 : entity xil_defaultlib.sysgen_abs_0161aa1824 
  port map (
    clr => '0',
    a => register7_q_net,
    clk => clk_net,
    ce => ce_net,
    op => absolute7_op_net
  );
end structural;
-- Generated from Simulink block PSB3_0/ov_detector_IFFT_im/Vector Absolute1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_absolute1 is
  port (
    d_1 : in std_logic_vector( 16-1 downto 0 );
    d_2 : in std_logic_vector( 16-1 downto 0 );
    d_3 : in std_logic_vector( 16-1 downto 0 );
    d_4 : in std_logic_vector( 16-1 downto 0 );
    d_5 : in std_logic_vector( 16-1 downto 0 );
    d_6 : in std_logic_vector( 16-1 downto 0 );
    d_7 : in std_logic_vector( 16-1 downto 0 );
    d_8 : in std_logic_vector( 16-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    q_1 : out std_logic_vector( 20-1 downto 0 );
    q_2 : out std_logic_vector( 20-1 downto 0 );
    q_3 : out std_logic_vector( 20-1 downto 0 );
    q_4 : out std_logic_vector( 20-1 downto 0 );
    q_5 : out std_logic_vector( 20-1 downto 0 );
    q_6 : out std_logic_vector( 20-1 downto 0 );
    q_7 : out std_logic_vector( 20-1 downto 0 );
    q_8 : out std_logic_vector( 20-1 downto 0 )
  );
end psb3_0_vector_absolute1;
architecture structural of psb3_0_vector_absolute1 is 
  signal mux4_y_net : std_logic_vector( 16-1 downto 0 );
  signal mux2_y_net : std_logic_vector( 16-1 downto 0 );
  signal mux5_y_net : std_logic_vector( 16-1 downto 0 );
  signal mux6_y_net : std_logic_vector( 16-1 downto 0 );
  signal mux7_y_net : std_logic_vector( 16-1 downto 0 );
  signal clk_net : std_logic;
  signal absolute4_op_net : std_logic_vector( 20-1 downto 0 );
  signal absolute7_op_net : std_logic_vector( 20-1 downto 0 );
  signal absolute5_op_net : std_logic_vector( 20-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 16-1 downto 0 );
  signal absolute0_op_net : std_logic_vector( 20-1 downto 0 );
  signal absolute6_op_net : std_logic_vector( 20-1 downto 0 );
  signal mux3_y_net : std_logic_vector( 16-1 downto 0 );
  signal absolute2_op_net : std_logic_vector( 20-1 downto 0 );
  signal absolute1_op_net : std_logic_vector( 20-1 downto 0 );
  signal absolute3_op_net : std_logic_vector( 20-1 downto 0 );
  signal mux0_y_net : std_logic_vector( 16-1 downto 0 );
  signal ce_net : std_logic;
begin
  q_1 <= absolute0_op_net;
  q_2 <= absolute1_op_net;
  q_3 <= absolute2_op_net;
  q_4 <= absolute3_op_net;
  q_5 <= absolute4_op_net;
  q_6 <= absolute5_op_net;
  q_7 <= absolute6_op_net;
  q_8 <= absolute7_op_net;
  mux0_y_net <= d_1;
  mux1_y_net <= d_2;
  mux2_y_net <= d_3;
  mux3_y_net <= d_4;
  mux4_y_net <= d_5;
  mux5_y_net <= d_6;
  mux6_y_net <= d_7;
  mux7_y_net <= d_8;
  clk_net <= clk_1;
  ce_net <= ce_1;
  absolute0 : entity xil_defaultlib.sysgen_abs_5e3e13aadc 
  port map (
    clr => '0',
    a => mux0_y_net,
    clk => clk_net,
    ce => ce_net,
    op => absolute0_op_net
  );
  absolute1 : entity xil_defaultlib.sysgen_abs_5e3e13aadc 
  port map (
    clr => '0',
    a => mux1_y_net,
    clk => clk_net,
    ce => ce_net,
    op => absolute1_op_net
  );
  absolute2 : entity xil_defaultlib.sysgen_abs_5e3e13aadc 
  port map (
    clr => '0',
    a => mux2_y_net,
    clk => clk_net,
    ce => ce_net,
    op => absolute2_op_net
  );
  absolute3 : entity xil_defaultlib.sysgen_abs_5e3e13aadc 
  port map (
    clr => '0',
    a => mux3_y_net,
    clk => clk_net,
    ce => ce_net,
    op => absolute3_op_net
  );
  absolute4 : entity xil_defaultlib.sysgen_abs_5e3e13aadc 
  port map (
    clr => '0',
    a => mux4_y_net,
    clk => clk_net,
    ce => ce_net,
    op => absolute4_op_net
  );
  absolute5 : entity xil_defaultlib.sysgen_abs_5e3e13aadc 
  port map (
    clr => '0',
    a => mux5_y_net,
    clk => clk_net,
    ce => ce_net,
    op => absolute5_op_net
  );
  absolute6 : entity xil_defaultlib.sysgen_abs_5e3e13aadc 
  port map (
    clr => '0',
    a => mux6_y_net,
    clk => clk_net,
    ce => ce_net,
    op => absolute6_op_net
  );
  absolute7 : entity xil_defaultlib.sysgen_abs_5e3e13aadc 
  port map (
    clr => '0',
    a => mux7_y_net,
    clk => clk_net,
    ce => ce_net,
    op => absolute7_op_net
  );
end structural;
-- Generated from Simulink block PSB3_0/ov_detector_IFFT_im/Vector Register
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_register is
  port (
    d_1 : in std_logic_vector( 20-1 downto 0 );
    rst : in std_logic_vector( 1-1 downto 0 );
    en : in std_logic;
    d_2 : in std_logic_vector( 20-1 downto 0 );
    d_3 : in std_logic_vector( 20-1 downto 0 );
    d_4 : in std_logic_vector( 20-1 downto 0 );
    d_5 : in std_logic_vector( 20-1 downto 0 );
    d_6 : in std_logic_vector( 20-1 downto 0 );
    d_7 : in std_logic_vector( 20-1 downto 0 );
    d_8 : in std_logic_vector( 20-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    q_1 : out std_logic_vector( 20-1 downto 0 );
    q_2 : out std_logic_vector( 20-1 downto 0 );
    q_3 : out std_logic_vector( 20-1 downto 0 );
    q_4 : out std_logic_vector( 20-1 downto 0 );
    q_5 : out std_logic_vector( 20-1 downto 0 );
    q_6 : out std_logic_vector( 20-1 downto 0 );
    q_7 : out std_logic_vector( 20-1 downto 0 );
    q_8 : out std_logic_vector( 20-1 downto 0 )
  );
end psb3_0_vector_register;
architecture structural of psb3_0_vector_register is 
  signal register7_q_net : std_logic_vector( 20-1 downto 0 );
  signal reinterpret16_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal register4_q_net : std_logic_vector( 20-1 downto 0 );
  signal register1_q_net : std_logic_vector( 20-1 downto 0 );
  signal gin_tl_reset_net : std_logic_vector( 1-1 downto 0 );
  signal test_systolicfft_vhdl_black_box_vo_net : std_logic;
  signal register2_q_net : std_logic_vector( 20-1 downto 0 );
  signal register5_q_net : std_logic_vector( 20-1 downto 0 );
  signal register6_q_net : std_logic_vector( 20-1 downto 0 );
  signal register3_q_net : std_logic_vector( 20-1 downto 0 );
  signal register0_q_net : std_logic_vector( 20-1 downto 0 );
  signal reinterpret21_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal reinterpret19_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal clk_net : std_logic;
  signal ce_net : std_logic;
  signal reinterpret17_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal reinterpret20_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal reinterpret22_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal reinterpret23_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal reinterpret18_output_port_net : std_logic_vector( 20-1 downto 0 );
begin
  q_1 <= register0_q_net;
  q_2 <= register1_q_net;
  q_3 <= register2_q_net;
  q_4 <= register3_q_net;
  q_5 <= register4_q_net;
  q_6 <= register5_q_net;
  q_7 <= register6_q_net;
  q_8 <= register7_q_net;
  reinterpret16_output_port_net <= d_1;
  gin_tl_reset_net <= rst;
  test_systolicfft_vhdl_black_box_vo_net <= en;
  reinterpret17_output_port_net <= d_2;
  reinterpret18_output_port_net <= d_3;
  reinterpret19_output_port_net <= d_4;
  reinterpret20_output_port_net <= d_5;
  reinterpret21_output_port_net <= d_6;
  reinterpret22_output_port_net <= d_7;
  reinterpret23_output_port_net <= d_8;
  clk_net <= clk_1;
  ce_net <= ce_1;
  register0 : entity xil_defaultlib.psb3_0_xlregister 
  generic map (
    d_width => 20,
    init_value => b"00000000000000000000"
  )
  port map (
    d => reinterpret16_output_port_net,
    rst => gin_tl_reset_net,
    en(0) => test_systolicfft_vhdl_black_box_vo_net,
    clk => clk_net,
    ce => ce_net,
    q => register0_q_net
  );
  register1 : entity xil_defaultlib.psb3_0_xlregister 
  generic map (
    d_width => 20,
    init_value => b"00000000000000000000"
  )
  port map (
    d => reinterpret17_output_port_net,
    rst => gin_tl_reset_net,
    en(0) => test_systolicfft_vhdl_black_box_vo_net,
    clk => clk_net,
    ce => ce_net,
    q => register1_q_net
  );
  register2 : entity xil_defaultlib.psb3_0_xlregister 
  generic map (
    d_width => 20,
    init_value => b"00000000000000000000"
  )
  port map (
    d => reinterpret18_output_port_net,
    rst => gin_tl_reset_net,
    en(0) => test_systolicfft_vhdl_black_box_vo_net,
    clk => clk_net,
    ce => ce_net,
    q => register2_q_net
  );
  register3 : entity xil_defaultlib.psb3_0_xlregister 
  generic map (
    d_width => 20,
    init_value => b"00000000000000000000"
  )
  port map (
    d => reinterpret19_output_port_net,
    rst => gin_tl_reset_net,
    en(0) => test_systolicfft_vhdl_black_box_vo_net,
    clk => clk_net,
    ce => ce_net,
    q => register3_q_net
  );
  register4 : entity xil_defaultlib.psb3_0_xlregister 
  generic map (
    d_width => 20,
    init_value => b"00000000000000000000"
  )
  port map (
    d => reinterpret20_output_port_net,
    rst => gin_tl_reset_net,
    en(0) => test_systolicfft_vhdl_black_box_vo_net,
    clk => clk_net,
    ce => ce_net,
    q => register4_q_net
  );
  register5 : entity xil_defaultlib.psb3_0_xlregister 
  generic map (
    d_width => 20,
    init_value => b"00000000000000000000"
  )
  port map (
    d => reinterpret21_output_port_net,
    rst => gin_tl_reset_net,
    en(0) => test_systolicfft_vhdl_black_box_vo_net,
    clk => clk_net,
    ce => ce_net,
    q => register5_q_net
  );
  register6 : entity xil_defaultlib.psb3_0_xlregister 
  generic map (
    d_width => 20,
    init_value => b"00000000000000000000"
  )
  port map (
    d => reinterpret22_output_port_net,
    rst => gin_tl_reset_net,
    en(0) => test_systolicfft_vhdl_black_box_vo_net,
    clk => clk_net,
    ce => ce_net,
    q => register6_q_net
  );
  register7 : entity xil_defaultlib.psb3_0_xlregister 
  generic map (
    d_width => 20,
    init_value => b"00000000000000000000"
  )
  port map (
    d => reinterpret23_output_port_net,
    rst => gin_tl_reset_net,
    en(0) => test_systolicfft_vhdl_black_box_vo_net,
    clk => clk_net,
    ce => ce_net,
    q => register7_q_net
  );
end structural;
-- Generated from Simulink block PSB3_0/ov_detector_IFFT_im/Vector Relational
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_relational is
  port (
    a_1 : in std_logic_vector( 20-1 downto 0 );
    b_1 : in std_logic_vector( 20-1 downto 0 );
    a_2 : in std_logic_vector( 20-1 downto 0 );
    a_3 : in std_logic_vector( 20-1 downto 0 );
    a_4 : in std_logic_vector( 20-1 downto 0 );
    a_5 : in std_logic_vector( 20-1 downto 0 );
    a_6 : in std_logic_vector( 20-1 downto 0 );
    a_7 : in std_logic_vector( 20-1 downto 0 );
    a_8 : in std_logic_vector( 20-1 downto 0 );
    b_2 : in std_logic_vector( 20-1 downto 0 );
    b_3 : in std_logic_vector( 20-1 downto 0 );
    b_4 : in std_logic_vector( 20-1 downto 0 );
    b_5 : in std_logic_vector( 20-1 downto 0 );
    b_6 : in std_logic_vector( 20-1 downto 0 );
    b_7 : in std_logic_vector( 20-1 downto 0 );
    b_8 : in std_logic_vector( 20-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    out_1 : out std_logic_vector( 1-1 downto 0 );
    out_2 : out std_logic_vector( 1-1 downto 0 );
    out_3 : out std_logic_vector( 1-1 downto 0 );
    out_4 : out std_logic_vector( 1-1 downto 0 );
    out_5 : out std_logic_vector( 1-1 downto 0 );
    out_6 : out std_logic_vector( 1-1 downto 0 );
    out_7 : out std_logic_vector( 1-1 downto 0 );
    out_8 : out std_logic_vector( 1-1 downto 0 )
  );
end psb3_0_vector_relational;
architecture structural of psb3_0_vector_relational is 
  signal absolute2_op_net : std_logic_vector( 20-1 downto 0 );
  signal relational5_op_net : std_logic_vector( 1-1 downto 0 );
  signal absolute2_op_net_x0 : std_logic_vector( 20-1 downto 0 );
  signal absolute7_op_net_x0 : std_logic_vector( 20-1 downto 0 );
  signal relational0_op_net : std_logic_vector( 1-1 downto 0 );
  signal absolute5_op_net_x0 : std_logic_vector( 20-1 downto 0 );
  signal absolute1_op_net : std_logic_vector( 20-1 downto 0 );
  signal absolute6_op_net : std_logic_vector( 20-1 downto 0 );
  signal relational2_op_net : std_logic_vector( 1-1 downto 0 );
  signal absolute3_op_net : std_logic_vector( 20-1 downto 0 );
  signal absolute1_op_net_x0 : std_logic_vector( 20-1 downto 0 );
  signal relational7_op_net : std_logic_vector( 1-1 downto 0 );
  signal absolute0_op_net : std_logic_vector( 20-1 downto 0 );
  signal absolute4_op_net : std_logic_vector( 20-1 downto 0 );
  signal absolute3_op_net_x0 : std_logic_vector( 20-1 downto 0 );
  signal absolute7_op_net : std_logic_vector( 20-1 downto 0 );
  signal clk_net : std_logic;
  signal ce_net : std_logic;
  signal relational1_op_net : std_logic_vector( 1-1 downto 0 );
  signal absolute0_op_net_x0 : std_logic_vector( 20-1 downto 0 );
  signal relational6_op_net : std_logic_vector( 1-1 downto 0 );
  signal absolute4_op_net_x0 : std_logic_vector( 20-1 downto 0 );
  signal absolute6_op_net_x0 : std_logic_vector( 20-1 downto 0 );
  signal relational3_op_net : std_logic_vector( 1-1 downto 0 );
  signal absolute5_op_net : std_logic_vector( 20-1 downto 0 );
  signal relational4_op_net : std_logic_vector( 1-1 downto 0 );
begin
  out_1 <= relational0_op_net;
  out_2 <= relational1_op_net;
  out_3 <= relational2_op_net;
  out_4 <= relational3_op_net;
  out_5 <= relational4_op_net;
  out_6 <= relational5_op_net;
  out_7 <= relational6_op_net;
  out_8 <= relational7_op_net;
  absolute0_op_net_x0 <= a_1;
  absolute0_op_net <= b_1;
  absolute1_op_net_x0 <= a_2;
  absolute2_op_net_x0 <= a_3;
  absolute3_op_net_x0 <= a_4;
  absolute4_op_net_x0 <= a_5;
  absolute5_op_net_x0 <= a_6;
  absolute6_op_net_x0 <= a_7;
  absolute7_op_net_x0 <= a_8;
  absolute1_op_net <= b_2;
  absolute2_op_net <= b_3;
  absolute3_op_net <= b_4;
  absolute4_op_net <= b_5;
  absolute5_op_net <= b_6;
  absolute6_op_net <= b_7;
  absolute7_op_net <= b_8;
  clk_net <= clk_1;
  ce_net <= ce_1;
  relational0 : entity xil_defaultlib.sysgen_relational_27302b866e 
  port map (
    clr => '0',
    a => absolute0_op_net_x0,
    b => absolute0_op_net,
    clk => clk_net,
    ce => ce_net,
    op => relational0_op_net
  );
  relational1 : entity xil_defaultlib.sysgen_relational_27302b866e 
  port map (
    clr => '0',
    a => absolute1_op_net_x0,
    b => absolute1_op_net,
    clk => clk_net,
    ce => ce_net,
    op => relational1_op_net
  );
  relational2 : entity xil_defaultlib.sysgen_relational_27302b866e 
  port map (
    clr => '0',
    a => absolute2_op_net_x0,
    b => absolute2_op_net,
    clk => clk_net,
    ce => ce_net,
    op => relational2_op_net
  );
  relational3 : entity xil_defaultlib.sysgen_relational_27302b866e 
  port map (
    clr => '0',
    a => absolute3_op_net_x0,
    b => absolute3_op_net,
    clk => clk_net,
    ce => ce_net,
    op => relational3_op_net
  );
  relational4 : entity xil_defaultlib.sysgen_relational_27302b866e 
  port map (
    clr => '0',
    a => absolute4_op_net_x0,
    b => absolute4_op_net,
    clk => clk_net,
    ce => ce_net,
    op => relational4_op_net
  );
  relational5 : entity xil_defaultlib.sysgen_relational_27302b866e 
  port map (
    clr => '0',
    a => absolute5_op_net_x0,
    b => absolute5_op_net,
    clk => clk_net,
    ce => ce_net,
    op => relational5_op_net
  );
  relational6 : entity xil_defaultlib.sysgen_relational_27302b866e 
  port map (
    clr => '0',
    a => absolute6_op_net_x0,
    b => absolute6_op_net,
    clk => clk_net,
    ce => ce_net,
    op => relational6_op_net
  );
  relational7 : entity xil_defaultlib.sysgen_relational_27302b866e 
  port map (
    clr => '0',
    a => absolute7_op_net_x0,
    b => absolute7_op_net,
    clk => clk_net,
    ce => ce_net,
    op => relational7_op_net
  );
end structural;
-- Generated from Simulink block PSB3_0/ov_detector_IFFT_im
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_ov_detector_ifft_im is
  port (
    rst : in std_logic_vector( 1-1 downto 0 );
    a_1 : in std_logic_vector( 20-1 downto 0 );
    b_1 : in std_logic_vector( 16-1 downto 0 );
    en : in std_logic;
    a_2 : in std_logic_vector( 20-1 downto 0 );
    a_3 : in std_logic_vector( 20-1 downto 0 );
    a_4 : in std_logic_vector( 20-1 downto 0 );
    a_5 : in std_logic_vector( 20-1 downto 0 );
    a_6 : in std_logic_vector( 20-1 downto 0 );
    a_7 : in std_logic_vector( 20-1 downto 0 );
    a_8 : in std_logic_vector( 20-1 downto 0 );
    b_2 : in std_logic_vector( 16-1 downto 0 );
    b_3 : in std_logic_vector( 16-1 downto 0 );
    b_4 : in std_logic_vector( 16-1 downto 0 );
    b_5 : in std_logic_vector( 16-1 downto 0 );
    b_6 : in std_logic_vector( 16-1 downto 0 );
    b_7 : in std_logic_vector( 16-1 downto 0 );
    b_8 : in std_logic_vector( 16-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    ov : out std_logic_vector( 1-1 downto 0 )
  );
end psb3_0_ov_detector_ifft_im;
architecture structural of psb3_0_ov_detector_ifft_im is 
  signal relational3_op_net : std_logic_vector( 1-1 downto 0 );
  signal constant17_op_net : std_logic_vector( 1-1 downto 0 );
  signal mux6_y_net : std_logic_vector( 16-1 downto 0 );
  signal mux7_y_net : std_logic_vector( 16-1 downto 0 );
  signal relational7_op_net : std_logic_vector( 1-1 downto 0 );
  signal mux5_y_net : std_logic_vector( 16-1 downto 0 );
  signal relational2_op_net : std_logic_vector( 1-1 downto 0 );
  signal mux3_y_net : std_logic_vector( 16-1 downto 0 );
  signal absolute5_op_net_x0 : std_logic_vector( 20-1 downto 0 );
  signal register7_q_net : std_logic_vector( 20-1 downto 0 );
  signal absolute4_op_net : std_logic_vector( 20-1 downto 0 );
  signal ce_net : std_logic;
  signal absolute7_op_net_x0 : std_logic_vector( 20-1 downto 0 );
  signal absolute3_op_net_x0 : std_logic_vector( 20-1 downto 0 );
  signal register1_q_net : std_logic_vector( 20-1 downto 0 );
  signal register5_q_net : std_logic_vector( 20-1 downto 0 );
  signal absolute4_op_net_x0 : std_logic_vector( 20-1 downto 0 );
  signal relational1_op_net : std_logic_vector( 1-1 downto 0 );
  signal register4_q_net : std_logic_vector( 20-1 downto 0 );
  signal relational4_op_net : std_logic_vector( 1-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 16-1 downto 0 );
  signal absolute5_op_net : std_logic_vector( 20-1 downto 0 );
  signal register0_q_net : std_logic_vector( 20-1 downto 0 );
  signal relational5_op_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret23_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal register6_q_net : std_logic_vector( 20-1 downto 0 );
  signal register3_q_net : std_logic_vector( 20-1 downto 0 );
  signal relational6_op_net : std_logic_vector( 1-1 downto 0 );
  signal absolute7_op_net : std_logic_vector( 20-1 downto 0 );
  signal register2_q_net : std_logic_vector( 20-1 downto 0 );
  signal absolute1_op_net : std_logic_vector( 20-1 downto 0 );
  signal mux4_y_net : std_logic_vector( 16-1 downto 0 );
  signal clk_net : std_logic;
  signal absolute0_op_net_x0 : std_logic_vector( 20-1 downto 0 );
  signal absolute2_op_net_x0 : std_logic_vector( 20-1 downto 0 );
  signal mux2_y_net : std_logic_vector( 16-1 downto 0 );
  signal absolute6_op_net_x0 : std_logic_vector( 20-1 downto 0 );
  signal absolute0_op_net : std_logic_vector( 20-1 downto 0 );
  signal absolute2_op_net : std_logic_vector( 20-1 downto 0 );
  signal absolute1_op_net_x0 : std_logic_vector( 20-1 downto 0 );
  signal absolute3_op_net : std_logic_vector( 20-1 downto 0 );
  signal absolute6_op_net : std_logic_vector( 20-1 downto 0 );
  signal relational0_op_net : std_logic_vector( 1-1 downto 0 );
  signal expression_dout_net : std_logic_vector( 1-1 downto 0 );
  signal gin_tl_reset_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret16_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal mux0_y_net : std_logic_vector( 16-1 downto 0 );
  signal test_systolicfft_vhdl_black_box_vo_net : std_logic;
  signal reinterpret17_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal reinterpret20_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal reinterpret19_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal reinterpret21_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal reinterpret22_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal reinterpret18_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal register_q_net : std_logic_vector( 1-1 downto 0 );
begin
  ov <= register_q_net;
  gin_tl_reset_net <= rst;
  reinterpret16_output_port_net <= a_1;
  mux0_y_net <= b_1;
  test_systolicfft_vhdl_black_box_vo_net <= en;
  reinterpret17_output_port_net <= a_2;
  reinterpret18_output_port_net <= a_3;
  reinterpret19_output_port_net <= a_4;
  reinterpret20_output_port_net <= a_5;
  reinterpret21_output_port_net <= a_6;
  reinterpret22_output_port_net <= a_7;
  reinterpret23_output_port_net <= a_8;
  mux1_y_net <= b_2;
  mux2_y_net <= b_3;
  mux3_y_net <= b_4;
  mux4_y_net <= b_5;
  mux5_y_net <= b_6;
  mux6_y_net <= b_7;
  mux7_y_net <= b_8;
  clk_net <= clk_1;
  ce_net <= ce_1;
  vector_absolute : entity xil_defaultlib.psb3_0_vector_absolute 
  port map (
    d_1 => register0_q_net,
    d_2 => register1_q_net,
    d_3 => register2_q_net,
    d_4 => register3_q_net,
    d_5 => register4_q_net,
    d_6 => register5_q_net,
    d_7 => register6_q_net,
    d_8 => register7_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    q_1 => absolute0_op_net_x0,
    q_2 => absolute1_op_net_x0,
    q_3 => absolute2_op_net_x0,
    q_4 => absolute3_op_net_x0,
    q_5 => absolute4_op_net_x0,
    q_6 => absolute5_op_net_x0,
    q_7 => absolute6_op_net_x0,
    q_8 => absolute7_op_net_x0
  );
  vector_absolute1 : entity xil_defaultlib.psb3_0_vector_absolute1 
  port map (
    d_1 => mux0_y_net,
    d_2 => mux1_y_net,
    d_3 => mux2_y_net,
    d_4 => mux3_y_net,
    d_5 => mux4_y_net,
    d_6 => mux5_y_net,
    d_7 => mux6_y_net,
    d_8 => mux7_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    q_1 => absolute0_op_net,
    q_2 => absolute1_op_net,
    q_3 => absolute2_op_net,
    q_4 => absolute3_op_net,
    q_5 => absolute4_op_net,
    q_6 => absolute5_op_net,
    q_7 => absolute6_op_net,
    q_8 => absolute7_op_net
  );
  vector_register : entity xil_defaultlib.psb3_0_vector_register 
  port map (
    d_1 => reinterpret16_output_port_net,
    rst => gin_tl_reset_net,
    en => test_systolicfft_vhdl_black_box_vo_net,
    d_2 => reinterpret17_output_port_net,
    d_3 => reinterpret18_output_port_net,
    d_4 => reinterpret19_output_port_net,
    d_5 => reinterpret20_output_port_net,
    d_6 => reinterpret21_output_port_net,
    d_7 => reinterpret22_output_port_net,
    d_8 => reinterpret23_output_port_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    q_1 => register0_q_net,
    q_2 => register1_q_net,
    q_3 => register2_q_net,
    q_4 => register3_q_net,
    q_5 => register4_q_net,
    q_6 => register5_q_net,
    q_7 => register6_q_net,
    q_8 => register7_q_net
  );
  vector_relational : entity xil_defaultlib.psb3_0_vector_relational 
  port map (
    a_1 => absolute0_op_net_x0,
    b_1 => absolute0_op_net,
    a_2 => absolute1_op_net_x0,
    a_3 => absolute2_op_net_x0,
    a_4 => absolute3_op_net_x0,
    a_5 => absolute4_op_net_x0,
    a_6 => absolute5_op_net_x0,
    a_7 => absolute6_op_net_x0,
    a_8 => absolute7_op_net_x0,
    b_2 => absolute1_op_net,
    b_3 => absolute2_op_net,
    b_4 => absolute3_op_net,
    b_5 => absolute4_op_net,
    b_6 => absolute5_op_net,
    b_7 => absolute6_op_net,
    b_8 => absolute7_op_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    out_1 => relational0_op_net,
    out_2 => relational1_op_net,
    out_3 => relational2_op_net,
    out_4 => relational3_op_net,
    out_5 => relational4_op_net,
    out_6 => relational5_op_net,
    out_7 => relational6_op_net,
    out_8 => relational7_op_net
  );
  constant17 : entity xil_defaultlib.sysgen_constant_71e89d757c 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant17_op_net
  );
  expression : entity xil_defaultlib.sysgen_expr_189d6fb430 
  port map (
    clr => '0',
    a1 => relational0_op_net,
    a2 => relational1_op_net,
    b1 => relational2_op_net,
    b2 => relational3_op_net,
    c1 => relational4_op_net,
    c2 => relational5_op_net,
    d1 => relational6_op_net,
    d2 => relational7_op_net,
    clk => clk_net,
    ce => ce_net,
    dout => expression_dout_net
  );
  register_x0 : entity xil_defaultlib.psb3_0_xlregister 
  generic map (
    d_width => 1,
    init_value => b"0"
  )
  port map (
    d => constant17_op_net,
    rst => gin_tl_reset_net,
    en => expression_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => register_q_net
  );
end structural;
-- Generated from Simulink block PSB3_0/ov_detector_IFFT_re/Vector Absolute
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_absolute_x0 is
  port (
    d_1 : in std_logic_vector( 20-1 downto 0 );
    d_2 : in std_logic_vector( 20-1 downto 0 );
    d_3 : in std_logic_vector( 20-1 downto 0 );
    d_4 : in std_logic_vector( 20-1 downto 0 );
    d_5 : in std_logic_vector( 20-1 downto 0 );
    d_6 : in std_logic_vector( 20-1 downto 0 );
    d_7 : in std_logic_vector( 20-1 downto 0 );
    d_8 : in std_logic_vector( 20-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    q_1 : out std_logic_vector( 20-1 downto 0 );
    q_2 : out std_logic_vector( 20-1 downto 0 );
    q_3 : out std_logic_vector( 20-1 downto 0 );
    q_4 : out std_logic_vector( 20-1 downto 0 );
    q_5 : out std_logic_vector( 20-1 downto 0 );
    q_6 : out std_logic_vector( 20-1 downto 0 );
    q_7 : out std_logic_vector( 20-1 downto 0 );
    q_8 : out std_logic_vector( 20-1 downto 0 )
  );
end psb3_0_vector_absolute_x0;
architecture structural of psb3_0_vector_absolute_x0 is 
  signal register3_q_net : std_logic_vector( 20-1 downto 0 );
  signal clk_net : std_logic;
  signal absolute0_op_net : std_logic_vector( 20-1 downto 0 );
  signal register4_q_net : std_logic_vector( 20-1 downto 0 );
  signal register7_q_net : std_logic_vector( 20-1 downto 0 );
  signal absolute4_op_net : std_logic_vector( 20-1 downto 0 );
  signal absolute1_op_net : std_logic_vector( 20-1 downto 0 );
  signal register2_q_net : std_logic_vector( 20-1 downto 0 );
  signal absolute3_op_net : std_logic_vector( 20-1 downto 0 );
  signal register1_q_net : std_logic_vector( 20-1 downto 0 );
  signal register5_q_net : std_logic_vector( 20-1 downto 0 );
  signal absolute5_op_net : std_logic_vector( 20-1 downto 0 );
  signal register6_q_net : std_logic_vector( 20-1 downto 0 );
  signal absolute6_op_net : std_logic_vector( 20-1 downto 0 );
  signal absolute2_op_net : std_logic_vector( 20-1 downto 0 );
  signal register0_q_net : std_logic_vector( 20-1 downto 0 );
  signal absolute7_op_net : std_logic_vector( 20-1 downto 0 );
  signal ce_net : std_logic;
begin
  q_1 <= absolute0_op_net;
  q_2 <= absolute1_op_net;
  q_3 <= absolute2_op_net;
  q_4 <= absolute3_op_net;
  q_5 <= absolute4_op_net;
  q_6 <= absolute5_op_net;
  q_7 <= absolute6_op_net;
  q_8 <= absolute7_op_net;
  register0_q_net <= d_1;
  register1_q_net <= d_2;
  register2_q_net <= d_3;
  register3_q_net <= d_4;
  register4_q_net <= d_5;
  register5_q_net <= d_6;
  register6_q_net <= d_7;
  register7_q_net <= d_8;
  clk_net <= clk_1;
  ce_net <= ce_1;
  absolute0 : entity xil_defaultlib.sysgen_abs_0161aa1824 
  port map (
    clr => '0',
    a => register0_q_net,
    clk => clk_net,
    ce => ce_net,
    op => absolute0_op_net
  );
  absolute1 : entity xil_defaultlib.sysgen_abs_0161aa1824 
  port map (
    clr => '0',
    a => register1_q_net,
    clk => clk_net,
    ce => ce_net,
    op => absolute1_op_net
  );
  absolute2 : entity xil_defaultlib.sysgen_abs_0161aa1824 
  port map (
    clr => '0',
    a => register2_q_net,
    clk => clk_net,
    ce => ce_net,
    op => absolute2_op_net
  );
  absolute3 : entity xil_defaultlib.sysgen_abs_0161aa1824 
  port map (
    clr => '0',
    a => register3_q_net,
    clk => clk_net,
    ce => ce_net,
    op => absolute3_op_net
  );
  absolute4 : entity xil_defaultlib.sysgen_abs_0161aa1824 
  port map (
    clr => '0',
    a => register4_q_net,
    clk => clk_net,
    ce => ce_net,
    op => absolute4_op_net
  );
  absolute5 : entity xil_defaultlib.sysgen_abs_0161aa1824 
  port map (
    clr => '0',
    a => register5_q_net,
    clk => clk_net,
    ce => ce_net,
    op => absolute5_op_net
  );
  absolute6 : entity xil_defaultlib.sysgen_abs_0161aa1824 
  port map (
    clr => '0',
    a => register6_q_net,
    clk => clk_net,
    ce => ce_net,
    op => absolute6_op_net
  );
  absolute7 : entity xil_defaultlib.sysgen_abs_0161aa1824 
  port map (
    clr => '0',
    a => register7_q_net,
    clk => clk_net,
    ce => ce_net,
    op => absolute7_op_net
  );
end structural;
-- Generated from Simulink block PSB3_0/ov_detector_IFFT_re/Vector Absolute1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_absolute1_x0 is
  port (
    d_1 : in std_logic_vector( 16-1 downto 0 );
    d_2 : in std_logic_vector( 16-1 downto 0 );
    d_3 : in std_logic_vector( 16-1 downto 0 );
    d_4 : in std_logic_vector( 16-1 downto 0 );
    d_5 : in std_logic_vector( 16-1 downto 0 );
    d_6 : in std_logic_vector( 16-1 downto 0 );
    d_7 : in std_logic_vector( 16-1 downto 0 );
    d_8 : in std_logic_vector( 16-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    q_1 : out std_logic_vector( 20-1 downto 0 );
    q_2 : out std_logic_vector( 20-1 downto 0 );
    q_3 : out std_logic_vector( 20-1 downto 0 );
    q_4 : out std_logic_vector( 20-1 downto 0 );
    q_5 : out std_logic_vector( 20-1 downto 0 );
    q_6 : out std_logic_vector( 20-1 downto 0 );
    q_7 : out std_logic_vector( 20-1 downto 0 );
    q_8 : out std_logic_vector( 20-1 downto 0 )
  );
end psb3_0_vector_absolute1_x0;
architecture structural of psb3_0_vector_absolute1_x0 is 
  signal ce_net : std_logic;
  signal mux2_y_net : std_logic_vector( 16-1 downto 0 );
  signal mux3_y_net : std_logic_vector( 16-1 downto 0 );
  signal mux5_y_net : std_logic_vector( 16-1 downto 0 );
  signal clk_net : std_logic;
  signal absolute4_op_net : std_logic_vector( 20-1 downto 0 );
  signal absolute2_op_net : std_logic_vector( 20-1 downto 0 );
  signal absolute5_op_net : std_logic_vector( 20-1 downto 0 );
  signal absolute1_op_net : std_logic_vector( 20-1 downto 0 );
  signal absolute6_op_net : std_logic_vector( 20-1 downto 0 );
  signal mux0_y_net : std_logic_vector( 16-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 16-1 downto 0 );
  signal mux4_y_net : std_logic_vector( 16-1 downto 0 );
  signal absolute7_op_net : std_logic_vector( 20-1 downto 0 );
  signal mux6_y_net : std_logic_vector( 16-1 downto 0 );
  signal absolute0_op_net : std_logic_vector( 20-1 downto 0 );
  signal absolute3_op_net : std_logic_vector( 20-1 downto 0 );
  signal mux7_y_net : std_logic_vector( 16-1 downto 0 );
begin
  q_1 <= absolute0_op_net;
  q_2 <= absolute1_op_net;
  q_3 <= absolute2_op_net;
  q_4 <= absolute3_op_net;
  q_5 <= absolute4_op_net;
  q_6 <= absolute5_op_net;
  q_7 <= absolute6_op_net;
  q_8 <= absolute7_op_net;
  mux0_y_net <= d_1;
  mux1_y_net <= d_2;
  mux2_y_net <= d_3;
  mux3_y_net <= d_4;
  mux4_y_net <= d_5;
  mux5_y_net <= d_6;
  mux6_y_net <= d_7;
  mux7_y_net <= d_8;
  clk_net <= clk_1;
  ce_net <= ce_1;
  absolute0 : entity xil_defaultlib.sysgen_abs_5e3e13aadc 
  port map (
    clr => '0',
    a => mux0_y_net,
    clk => clk_net,
    ce => ce_net,
    op => absolute0_op_net
  );
  absolute1 : entity xil_defaultlib.sysgen_abs_5e3e13aadc 
  port map (
    clr => '0',
    a => mux1_y_net,
    clk => clk_net,
    ce => ce_net,
    op => absolute1_op_net
  );
  absolute2 : entity xil_defaultlib.sysgen_abs_5e3e13aadc 
  port map (
    clr => '0',
    a => mux2_y_net,
    clk => clk_net,
    ce => ce_net,
    op => absolute2_op_net
  );
  absolute3 : entity xil_defaultlib.sysgen_abs_5e3e13aadc 
  port map (
    clr => '0',
    a => mux3_y_net,
    clk => clk_net,
    ce => ce_net,
    op => absolute3_op_net
  );
  absolute4 : entity xil_defaultlib.sysgen_abs_5e3e13aadc 
  port map (
    clr => '0',
    a => mux4_y_net,
    clk => clk_net,
    ce => ce_net,
    op => absolute4_op_net
  );
  absolute5 : entity xil_defaultlib.sysgen_abs_5e3e13aadc 
  port map (
    clr => '0',
    a => mux5_y_net,
    clk => clk_net,
    ce => ce_net,
    op => absolute5_op_net
  );
  absolute6 : entity xil_defaultlib.sysgen_abs_5e3e13aadc 
  port map (
    clr => '0',
    a => mux6_y_net,
    clk => clk_net,
    ce => ce_net,
    op => absolute6_op_net
  );
  absolute7 : entity xil_defaultlib.sysgen_abs_5e3e13aadc 
  port map (
    clr => '0',
    a => mux7_y_net,
    clk => clk_net,
    ce => ce_net,
    op => absolute7_op_net
  );
end structural;
-- Generated from Simulink block PSB3_0/ov_detector_IFFT_re/Vector Register
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_register_x0 is
  port (
    d_1 : in std_logic_vector( 20-1 downto 0 );
    rst : in std_logic_vector( 1-1 downto 0 );
    en : in std_logic;
    d_2 : in std_logic_vector( 20-1 downto 0 );
    d_3 : in std_logic_vector( 20-1 downto 0 );
    d_4 : in std_logic_vector( 20-1 downto 0 );
    d_5 : in std_logic_vector( 20-1 downto 0 );
    d_6 : in std_logic_vector( 20-1 downto 0 );
    d_7 : in std_logic_vector( 20-1 downto 0 );
    d_8 : in std_logic_vector( 20-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    q_1 : out std_logic_vector( 20-1 downto 0 );
    q_2 : out std_logic_vector( 20-1 downto 0 );
    q_3 : out std_logic_vector( 20-1 downto 0 );
    q_4 : out std_logic_vector( 20-1 downto 0 );
    q_5 : out std_logic_vector( 20-1 downto 0 );
    q_6 : out std_logic_vector( 20-1 downto 0 );
    q_7 : out std_logic_vector( 20-1 downto 0 );
    q_8 : out std_logic_vector( 20-1 downto 0 )
  );
end psb3_0_vector_register_x0;
architecture structural of psb3_0_vector_register_x0 is 
  signal register6_q_net : std_logic_vector( 20-1 downto 0 );
  signal register7_q_net : std_logic_vector( 20-1 downto 0 );
  signal reinterpret24_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal gin_tl_reset_net : std_logic_vector( 1-1 downto 0 );
  signal test_systolicfft_vhdl_black_box_vo_net : std_logic;
  signal reinterpret25_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal register0_q_net : std_logic_vector( 20-1 downto 0 );
  signal register1_q_net : std_logic_vector( 20-1 downto 0 );
  signal register2_q_net : std_logic_vector( 20-1 downto 0 );
  signal register3_q_net : std_logic_vector( 20-1 downto 0 );
  signal register4_q_net : std_logic_vector( 20-1 downto 0 );
  signal register5_q_net : std_logic_vector( 20-1 downto 0 );
  signal reinterpret30_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal reinterpret29_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal ce_net : std_logic;
  signal clk_net : std_logic;
  signal reinterpret28_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal reinterpret27_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal reinterpret31_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal reinterpret26_output_port_net : std_logic_vector( 20-1 downto 0 );
begin
  q_1 <= register0_q_net;
  q_2 <= register1_q_net;
  q_3 <= register2_q_net;
  q_4 <= register3_q_net;
  q_5 <= register4_q_net;
  q_6 <= register5_q_net;
  q_7 <= register6_q_net;
  q_8 <= register7_q_net;
  reinterpret24_output_port_net <= d_1;
  gin_tl_reset_net <= rst;
  test_systolicfft_vhdl_black_box_vo_net <= en;
  reinterpret25_output_port_net <= d_2;
  reinterpret26_output_port_net <= d_3;
  reinterpret27_output_port_net <= d_4;
  reinterpret28_output_port_net <= d_5;
  reinterpret29_output_port_net <= d_6;
  reinterpret30_output_port_net <= d_7;
  reinterpret31_output_port_net <= d_8;
  clk_net <= clk_1;
  ce_net <= ce_1;
  register0 : entity xil_defaultlib.psb3_0_xlregister 
  generic map (
    d_width => 20,
    init_value => b"00000000000000000000"
  )
  port map (
    d => reinterpret24_output_port_net,
    rst => gin_tl_reset_net,
    en(0) => test_systolicfft_vhdl_black_box_vo_net,
    clk => clk_net,
    ce => ce_net,
    q => register0_q_net
  );
  register1 : entity xil_defaultlib.psb3_0_xlregister 
  generic map (
    d_width => 20,
    init_value => b"00000000000000000000"
  )
  port map (
    d => reinterpret25_output_port_net,
    rst => gin_tl_reset_net,
    en(0) => test_systolicfft_vhdl_black_box_vo_net,
    clk => clk_net,
    ce => ce_net,
    q => register1_q_net
  );
  register2 : entity xil_defaultlib.psb3_0_xlregister 
  generic map (
    d_width => 20,
    init_value => b"00000000000000000000"
  )
  port map (
    d => reinterpret26_output_port_net,
    rst => gin_tl_reset_net,
    en(0) => test_systolicfft_vhdl_black_box_vo_net,
    clk => clk_net,
    ce => ce_net,
    q => register2_q_net
  );
  register3 : entity xil_defaultlib.psb3_0_xlregister 
  generic map (
    d_width => 20,
    init_value => b"00000000000000000000"
  )
  port map (
    d => reinterpret27_output_port_net,
    rst => gin_tl_reset_net,
    en(0) => test_systolicfft_vhdl_black_box_vo_net,
    clk => clk_net,
    ce => ce_net,
    q => register3_q_net
  );
  register4 : entity xil_defaultlib.psb3_0_xlregister 
  generic map (
    d_width => 20,
    init_value => b"00000000000000000000"
  )
  port map (
    d => reinterpret28_output_port_net,
    rst => gin_tl_reset_net,
    en(0) => test_systolicfft_vhdl_black_box_vo_net,
    clk => clk_net,
    ce => ce_net,
    q => register4_q_net
  );
  register5 : entity xil_defaultlib.psb3_0_xlregister 
  generic map (
    d_width => 20,
    init_value => b"00000000000000000000"
  )
  port map (
    d => reinterpret29_output_port_net,
    rst => gin_tl_reset_net,
    en(0) => test_systolicfft_vhdl_black_box_vo_net,
    clk => clk_net,
    ce => ce_net,
    q => register5_q_net
  );
  register6 : entity xil_defaultlib.psb3_0_xlregister 
  generic map (
    d_width => 20,
    init_value => b"00000000000000000000"
  )
  port map (
    d => reinterpret30_output_port_net,
    rst => gin_tl_reset_net,
    en(0) => test_systolicfft_vhdl_black_box_vo_net,
    clk => clk_net,
    ce => ce_net,
    q => register6_q_net
  );
  register7 : entity xil_defaultlib.psb3_0_xlregister 
  generic map (
    d_width => 20,
    init_value => b"00000000000000000000"
  )
  port map (
    d => reinterpret31_output_port_net,
    rst => gin_tl_reset_net,
    en(0) => test_systolicfft_vhdl_black_box_vo_net,
    clk => clk_net,
    ce => ce_net,
    q => register7_q_net
  );
end structural;
-- Generated from Simulink block PSB3_0/ov_detector_IFFT_re/Vector Relational
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_relational_x0 is
  port (
    a_1 : in std_logic_vector( 20-1 downto 0 );
    b_1 : in std_logic_vector( 20-1 downto 0 );
    a_2 : in std_logic_vector( 20-1 downto 0 );
    a_3 : in std_logic_vector( 20-1 downto 0 );
    a_4 : in std_logic_vector( 20-1 downto 0 );
    a_5 : in std_logic_vector( 20-1 downto 0 );
    a_6 : in std_logic_vector( 20-1 downto 0 );
    a_7 : in std_logic_vector( 20-1 downto 0 );
    a_8 : in std_logic_vector( 20-1 downto 0 );
    b_2 : in std_logic_vector( 20-1 downto 0 );
    b_3 : in std_logic_vector( 20-1 downto 0 );
    b_4 : in std_logic_vector( 20-1 downto 0 );
    b_5 : in std_logic_vector( 20-1 downto 0 );
    b_6 : in std_logic_vector( 20-1 downto 0 );
    b_7 : in std_logic_vector( 20-1 downto 0 );
    b_8 : in std_logic_vector( 20-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    out_1 : out std_logic_vector( 1-1 downto 0 );
    out_2 : out std_logic_vector( 1-1 downto 0 );
    out_3 : out std_logic_vector( 1-1 downto 0 );
    out_4 : out std_logic_vector( 1-1 downto 0 );
    out_5 : out std_logic_vector( 1-1 downto 0 );
    out_6 : out std_logic_vector( 1-1 downto 0 );
    out_7 : out std_logic_vector( 1-1 downto 0 );
    out_8 : out std_logic_vector( 1-1 downto 0 )
  );
end psb3_0_vector_relational_x0;
architecture structural of psb3_0_vector_relational_x0 is 
  signal absolute1_op_net : std_logic_vector( 20-1 downto 0 );
  signal absolute2_op_net : std_logic_vector( 20-1 downto 0 );
  signal relational6_op_net : std_logic_vector( 1-1 downto 0 );
  signal relational3_op_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal relational2_op_net : std_logic_vector( 1-1 downto 0 );
  signal absolute3_op_net : std_logic_vector( 20-1 downto 0 );
  signal relational7_op_net : std_logic_vector( 1-1 downto 0 );
  signal absolute4_op_net_x0 : std_logic_vector( 20-1 downto 0 );
  signal ce_net : std_logic;
  signal absolute0_op_net : std_logic_vector( 20-1 downto 0 );
  signal absolute5_op_net : std_logic_vector( 20-1 downto 0 );
  signal absolute5_op_net_x0 : std_logic_vector( 20-1 downto 0 );
  signal relational0_op_net : std_logic_vector( 1-1 downto 0 );
  signal relational1_op_net : std_logic_vector( 1-1 downto 0 );
  signal absolute6_op_net_x0 : std_logic_vector( 20-1 downto 0 );
  signal absolute0_op_net_x0 : std_logic_vector( 20-1 downto 0 );
  signal absolute4_op_net : std_logic_vector( 20-1 downto 0 );
  signal absolute6_op_net : std_logic_vector( 20-1 downto 0 );
  signal absolute7_op_net : std_logic_vector( 20-1 downto 0 );
  signal relational5_op_net : std_logic_vector( 1-1 downto 0 );
  signal absolute7_op_net_x0 : std_logic_vector( 20-1 downto 0 );
  signal absolute2_op_net_x0 : std_logic_vector( 20-1 downto 0 );
  signal absolute3_op_net_x0 : std_logic_vector( 20-1 downto 0 );
  signal absolute1_op_net_x0 : std_logic_vector( 20-1 downto 0 );
  signal relational4_op_net : std_logic_vector( 1-1 downto 0 );
begin
  out_1 <= relational0_op_net;
  out_2 <= relational1_op_net;
  out_3 <= relational2_op_net;
  out_4 <= relational3_op_net;
  out_5 <= relational4_op_net;
  out_6 <= relational5_op_net;
  out_7 <= relational6_op_net;
  out_8 <= relational7_op_net;
  absolute0_op_net_x0 <= a_1;
  absolute0_op_net <= b_1;
  absolute1_op_net_x0 <= a_2;
  absolute2_op_net_x0 <= a_3;
  absolute3_op_net_x0 <= a_4;
  absolute4_op_net_x0 <= a_5;
  absolute5_op_net_x0 <= a_6;
  absolute6_op_net_x0 <= a_7;
  absolute7_op_net_x0 <= a_8;
  absolute1_op_net <= b_2;
  absolute2_op_net <= b_3;
  absolute3_op_net <= b_4;
  absolute4_op_net <= b_5;
  absolute5_op_net <= b_6;
  absolute6_op_net <= b_7;
  absolute7_op_net <= b_8;
  clk_net <= clk_1;
  ce_net <= ce_1;
  relational0 : entity xil_defaultlib.sysgen_relational_27302b866e 
  port map (
    clr => '0',
    a => absolute0_op_net_x0,
    b => absolute0_op_net,
    clk => clk_net,
    ce => ce_net,
    op => relational0_op_net
  );
  relational1 : entity xil_defaultlib.sysgen_relational_27302b866e 
  port map (
    clr => '0',
    a => absolute1_op_net_x0,
    b => absolute1_op_net,
    clk => clk_net,
    ce => ce_net,
    op => relational1_op_net
  );
  relational2 : entity xil_defaultlib.sysgen_relational_27302b866e 
  port map (
    clr => '0',
    a => absolute2_op_net_x0,
    b => absolute2_op_net,
    clk => clk_net,
    ce => ce_net,
    op => relational2_op_net
  );
  relational3 : entity xil_defaultlib.sysgen_relational_27302b866e 
  port map (
    clr => '0',
    a => absolute3_op_net_x0,
    b => absolute3_op_net,
    clk => clk_net,
    ce => ce_net,
    op => relational3_op_net
  );
  relational4 : entity xil_defaultlib.sysgen_relational_27302b866e 
  port map (
    clr => '0',
    a => absolute4_op_net_x0,
    b => absolute4_op_net,
    clk => clk_net,
    ce => ce_net,
    op => relational4_op_net
  );
  relational5 : entity xil_defaultlib.sysgen_relational_27302b866e 
  port map (
    clr => '0',
    a => absolute5_op_net_x0,
    b => absolute5_op_net,
    clk => clk_net,
    ce => ce_net,
    op => relational5_op_net
  );
  relational6 : entity xil_defaultlib.sysgen_relational_27302b866e 
  port map (
    clr => '0',
    a => absolute6_op_net_x0,
    b => absolute6_op_net,
    clk => clk_net,
    ce => ce_net,
    op => relational6_op_net
  );
  relational7 : entity xil_defaultlib.sysgen_relational_27302b866e 
  port map (
    clr => '0',
    a => absolute7_op_net_x0,
    b => absolute7_op_net,
    clk => clk_net,
    ce => ce_net,
    op => relational7_op_net
  );
end structural;
-- Generated from Simulink block PSB3_0/ov_detector_IFFT_re
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_ov_detector_ifft_re is
  port (
    rst : in std_logic_vector( 1-1 downto 0 );
    a_1 : in std_logic_vector( 20-1 downto 0 );
    b_1 : in std_logic_vector( 16-1 downto 0 );
    en : in std_logic;
    a_2 : in std_logic_vector( 20-1 downto 0 );
    a_3 : in std_logic_vector( 20-1 downto 0 );
    a_4 : in std_logic_vector( 20-1 downto 0 );
    a_5 : in std_logic_vector( 20-1 downto 0 );
    a_6 : in std_logic_vector( 20-1 downto 0 );
    a_7 : in std_logic_vector( 20-1 downto 0 );
    a_8 : in std_logic_vector( 20-1 downto 0 );
    b_2 : in std_logic_vector( 16-1 downto 0 );
    b_3 : in std_logic_vector( 16-1 downto 0 );
    b_4 : in std_logic_vector( 16-1 downto 0 );
    b_5 : in std_logic_vector( 16-1 downto 0 );
    b_6 : in std_logic_vector( 16-1 downto 0 );
    b_7 : in std_logic_vector( 16-1 downto 0 );
    b_8 : in std_logic_vector( 16-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    ov : out std_logic_vector( 1-1 downto 0 )
  );
end psb3_0_ov_detector_ifft_re;
architecture structural of psb3_0_ov_detector_ifft_re is 
  signal mux1_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret31_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal mux0_y_net : std_logic_vector( 16-1 downto 0 );
  signal register_q_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret24_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal test_systolicfft_vhdl_black_box_vo_net : std_logic;
  signal reinterpret25_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal reinterpret26_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal reinterpret27_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal reinterpret28_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal reinterpret29_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal gin_tl_reset_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret30_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal absolute0_op_net : std_logic_vector( 20-1 downto 0 );
  signal mux2_y_net : std_logic_vector( 16-1 downto 0 );
  signal absolute6_op_net : std_logic_vector( 20-1 downto 0 );
  signal mux6_y_net : std_logic_vector( 16-1 downto 0 );
  signal absolute1_op_net_x0 : std_logic_vector( 20-1 downto 0 );
  signal register3_q_net : std_logic_vector( 20-1 downto 0 );
  signal absolute3_op_net : std_logic_vector( 20-1 downto 0 );
  signal relational5_op_net : std_logic_vector( 1-1 downto 0 );
  signal relational6_op_net : std_logic_vector( 1-1 downto 0 );
  signal absolute1_op_net : std_logic_vector( 20-1 downto 0 );
  signal mux7_y_net : std_logic_vector( 16-1 downto 0 );
  signal register2_q_net : std_logic_vector( 20-1 downto 0 );
  signal absolute7_op_net : std_logic_vector( 20-1 downto 0 );
  signal relational4_op_net : std_logic_vector( 1-1 downto 0 );
  signal register1_q_net : std_logic_vector( 20-1 downto 0 );
  signal clk_net : std_logic;
  signal absolute0_op_net_x0 : std_logic_vector( 20-1 downto 0 );
  signal register0_q_net : std_logic_vector( 20-1 downto 0 );
  signal register6_q_net : std_logic_vector( 20-1 downto 0 );
  signal absolute2_op_net : std_logic_vector( 20-1 downto 0 );
  signal relational0_op_net : std_logic_vector( 1-1 downto 0 );
  signal relational2_op_net : std_logic_vector( 1-1 downto 0 );
  signal absolute5_op_net_x0 : std_logic_vector( 20-1 downto 0 );
  signal register7_q_net : std_logic_vector( 20-1 downto 0 );
  signal absolute2_op_net_x0 : std_logic_vector( 20-1 downto 0 );
  signal absolute4_op_net : std_logic_vector( 20-1 downto 0 );
  signal register4_q_net : std_logic_vector( 20-1 downto 0 );
  signal mux4_y_net : std_logic_vector( 16-1 downto 0 );
  signal mux3_y_net : std_logic_vector( 16-1 downto 0 );
  signal mux5_y_net : std_logic_vector( 16-1 downto 0 );
  signal relational1_op_net : std_logic_vector( 1-1 downto 0 );
  signal absolute7_op_net_x0 : std_logic_vector( 20-1 downto 0 );
  signal relational3_op_net : std_logic_vector( 1-1 downto 0 );
  signal relational7_op_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal register5_q_net : std_logic_vector( 20-1 downto 0 );
  signal constant17_op_net : std_logic_vector( 1-1 downto 0 );
  signal absolute5_op_net : std_logic_vector( 20-1 downto 0 );
  signal absolute6_op_net_x0 : std_logic_vector( 20-1 downto 0 );
  signal absolute3_op_net_x0 : std_logic_vector( 20-1 downto 0 );
  signal absolute4_op_net_x0 : std_logic_vector( 20-1 downto 0 );
  signal expression_dout_net : std_logic_vector( 1-1 downto 0 );
begin
  ov <= register_q_net;
  gin_tl_reset_net <= rst;
  reinterpret24_output_port_net <= a_1;
  mux0_y_net <= b_1;
  test_systolicfft_vhdl_black_box_vo_net <= en;
  reinterpret25_output_port_net <= a_2;
  reinterpret26_output_port_net <= a_3;
  reinterpret27_output_port_net <= a_4;
  reinterpret28_output_port_net <= a_5;
  reinterpret29_output_port_net <= a_6;
  reinterpret30_output_port_net <= a_7;
  reinterpret31_output_port_net <= a_8;
  mux1_y_net <= b_2;
  mux2_y_net <= b_3;
  mux3_y_net <= b_4;
  mux4_y_net <= b_5;
  mux5_y_net <= b_6;
  mux6_y_net <= b_7;
  mux7_y_net <= b_8;
  clk_net <= clk_1;
  ce_net <= ce_1;
  vector_absolute : entity xil_defaultlib.psb3_0_vector_absolute_x0 
  port map (
    d_1 => register0_q_net,
    d_2 => register1_q_net,
    d_3 => register2_q_net,
    d_4 => register3_q_net,
    d_5 => register4_q_net,
    d_6 => register5_q_net,
    d_7 => register6_q_net,
    d_8 => register7_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    q_1 => absolute0_op_net_x0,
    q_2 => absolute1_op_net_x0,
    q_3 => absolute2_op_net_x0,
    q_4 => absolute3_op_net_x0,
    q_5 => absolute4_op_net_x0,
    q_6 => absolute5_op_net_x0,
    q_7 => absolute6_op_net_x0,
    q_8 => absolute7_op_net_x0
  );
  vector_absolute1 : entity xil_defaultlib.psb3_0_vector_absolute1_x0 
  port map (
    d_1 => mux0_y_net,
    d_2 => mux1_y_net,
    d_3 => mux2_y_net,
    d_4 => mux3_y_net,
    d_5 => mux4_y_net,
    d_6 => mux5_y_net,
    d_7 => mux6_y_net,
    d_8 => mux7_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    q_1 => absolute0_op_net,
    q_2 => absolute1_op_net,
    q_3 => absolute2_op_net,
    q_4 => absolute3_op_net,
    q_5 => absolute4_op_net,
    q_6 => absolute5_op_net,
    q_7 => absolute6_op_net,
    q_8 => absolute7_op_net
  );
  vector_register : entity xil_defaultlib.psb3_0_vector_register_x0 
  port map (
    d_1 => reinterpret24_output_port_net,
    rst => gin_tl_reset_net,
    en => test_systolicfft_vhdl_black_box_vo_net,
    d_2 => reinterpret25_output_port_net,
    d_3 => reinterpret26_output_port_net,
    d_4 => reinterpret27_output_port_net,
    d_5 => reinterpret28_output_port_net,
    d_6 => reinterpret29_output_port_net,
    d_7 => reinterpret30_output_port_net,
    d_8 => reinterpret31_output_port_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    q_1 => register0_q_net,
    q_2 => register1_q_net,
    q_3 => register2_q_net,
    q_4 => register3_q_net,
    q_5 => register4_q_net,
    q_6 => register5_q_net,
    q_7 => register6_q_net,
    q_8 => register7_q_net
  );
  vector_relational : entity xil_defaultlib.psb3_0_vector_relational_x0 
  port map (
    a_1 => absolute0_op_net_x0,
    b_1 => absolute0_op_net,
    a_2 => absolute1_op_net_x0,
    a_3 => absolute2_op_net_x0,
    a_4 => absolute3_op_net_x0,
    a_5 => absolute4_op_net_x0,
    a_6 => absolute5_op_net_x0,
    a_7 => absolute6_op_net_x0,
    a_8 => absolute7_op_net_x0,
    b_2 => absolute1_op_net,
    b_3 => absolute2_op_net,
    b_4 => absolute3_op_net,
    b_5 => absolute4_op_net,
    b_6 => absolute5_op_net,
    b_7 => absolute6_op_net,
    b_8 => absolute7_op_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    out_1 => relational0_op_net,
    out_2 => relational1_op_net,
    out_3 => relational2_op_net,
    out_4 => relational3_op_net,
    out_5 => relational4_op_net,
    out_6 => relational5_op_net,
    out_7 => relational6_op_net,
    out_8 => relational7_op_net
  );
  constant17 : entity xil_defaultlib.sysgen_constant_71e89d757c 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant17_op_net
  );
  expression : entity xil_defaultlib.sysgen_expr_189d6fb430 
  port map (
    clr => '0',
    a1 => relational0_op_net,
    a2 => relational1_op_net,
    b1 => relational2_op_net,
    b2 => relational3_op_net,
    c1 => relational4_op_net,
    c2 => relational5_op_net,
    d1 => relational6_op_net,
    d2 => relational7_op_net,
    clk => clk_net,
    ce => ce_net,
    dout => expression_dout_net
  );
  register_x0 : entity xil_defaultlib.psb3_0_xlregister 
  generic map (
    d_width => 1,
    init_value => b"0"
  )
  port map (
    d => constant17_op_net,
    rst => gin_tl_reset_net,
    en => expression_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => register_q_net
  );
end structural;
-- Generated from Simulink block PSB3_0/reordering extending buffer imag_1/Scalar to Vector4
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_scalar_to_vector4_x0 is
  port (
    i : in std_logic_vector( 256-1 downto 0 );
    o_1 : out std_logic_vector( 16-1 downto 0 );
    o_2 : out std_logic_vector( 16-1 downto 0 );
    o_3 : out std_logic_vector( 16-1 downto 0 );
    o_4 : out std_logic_vector( 16-1 downto 0 );
    o_5 : out std_logic_vector( 16-1 downto 0 );
    o_6 : out std_logic_vector( 16-1 downto 0 );
    o_7 : out std_logic_vector( 16-1 downto 0 );
    o_8 : out std_logic_vector( 16-1 downto 0 );
    o_9 : out std_logic_vector( 16-1 downto 0 );
    o_10 : out std_logic_vector( 16-1 downto 0 );
    o_11 : out std_logic_vector( 16-1 downto 0 );
    o_12 : out std_logic_vector( 16-1 downto 0 );
    o_13 : out std_logic_vector( 16-1 downto 0 );
    o_14 : out std_logic_vector( 16-1 downto 0 );
    o_15 : out std_logic_vector( 16-1 downto 0 );
    o_16 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_scalar_to_vector4_x0;
architecture structural of psb3_0_scalar_to_vector4_x0 is 
  signal slice4_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 16-1 downto 0 );
  signal mux5_y_net : std_logic_vector( 256-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 16-1 downto 0 );
begin
  o_1 <= slice0_y_net;
  o_2 <= slice1_y_net;
  o_3 <= slice2_y_net;
  o_4 <= slice3_y_net;
  o_5 <= slice4_y_net;
  o_6 <= slice5_y_net;
  o_7 <= slice6_y_net;
  o_8 <= slice7_y_net;
  o_9 <= slice8_y_net;
  o_10 <= slice9_y_net;
  o_11 <= slice10_y_net;
  o_12 <= slice11_y_net;
  o_13 <= slice12_y_net;
  o_14 <= slice13_y_net;
  o_15 <= slice14_y_net;
  o_16 <= slice15_y_net;
  mux5_y_net <= i;
  slice0 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 15,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice0_y_net
  );
  slice1 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 16,
    new_msb => 31,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice1_y_net
  );
  slice2 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 32,
    new_msb => 47,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice2_y_net
  );
  slice3 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 48,
    new_msb => 63,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice3_y_net
  );
  slice4 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 64,
    new_msb => 79,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice4_y_net
  );
  slice5 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 80,
    new_msb => 95,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice5_y_net
  );
  slice6 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 96,
    new_msb => 111,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice6_y_net
  );
  slice7 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 112,
    new_msb => 127,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice7_y_net
  );
  slice8 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 128,
    new_msb => 143,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice8_y_net
  );
  slice9 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 144,
    new_msb => 159,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice9_y_net
  );
  slice10 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 160,
    new_msb => 175,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice10_y_net
  );
  slice11 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 176,
    new_msb => 191,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice11_y_net
  );
  slice12 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 192,
    new_msb => 207,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice12_y_net
  );
  slice13 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 208,
    new_msb => 223,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice13_y_net
  );
  slice14 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 224,
    new_msb => 239,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice14_y_net
  );
  slice15 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 240,
    new_msb => 255,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice15_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/reordering extending buffer imag_1/Vector Reinterpret
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_reinterpret_x3 is
  port (
    in_1 : in std_logic_vector( 16-1 downto 0 );
    in_2 : in std_logic_vector( 16-1 downto 0 );
    in_3 : in std_logic_vector( 16-1 downto 0 );
    in_4 : in std_logic_vector( 16-1 downto 0 );
    in_5 : in std_logic_vector( 16-1 downto 0 );
    in_6 : in std_logic_vector( 16-1 downto 0 );
    in_7 : in std_logic_vector( 16-1 downto 0 );
    in_8 : in std_logic_vector( 16-1 downto 0 );
    in_9 : in std_logic_vector( 16-1 downto 0 );
    in_10 : in std_logic_vector( 16-1 downto 0 );
    in_11 : in std_logic_vector( 16-1 downto 0 );
    in_12 : in std_logic_vector( 16-1 downto 0 );
    in_13 : in std_logic_vector( 16-1 downto 0 );
    in_14 : in std_logic_vector( 16-1 downto 0 );
    in_15 : in std_logic_vector( 16-1 downto 0 );
    in_16 : in std_logic_vector( 16-1 downto 0 );
    out_1 : out std_logic_vector( 16-1 downto 0 );
    out_2 : out std_logic_vector( 16-1 downto 0 );
    out_3 : out std_logic_vector( 16-1 downto 0 );
    out_4 : out std_logic_vector( 16-1 downto 0 );
    out_5 : out std_logic_vector( 16-1 downto 0 );
    out_6 : out std_logic_vector( 16-1 downto 0 );
    out_7 : out std_logic_vector( 16-1 downto 0 );
    out_8 : out std_logic_vector( 16-1 downto 0 );
    out_9 : out std_logic_vector( 16-1 downto 0 );
    out_10 : out std_logic_vector( 16-1 downto 0 );
    out_11 : out std_logic_vector( 16-1 downto 0 );
    out_12 : out std_logic_vector( 16-1 downto 0 );
    out_13 : out std_logic_vector( 16-1 downto 0 );
    out_14 : out std_logic_vector( 16-1 downto 0 );
    out_15 : out std_logic_vector( 16-1 downto 0 );
    out_16 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_vector_reinterpret_x3;
architecture structural of psb3_0_vector_reinterpret_x3 is 
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 16-1 downto 0 );
begin
  out_1 <= reinterpret0_output_port_net;
  out_2 <= reinterpret1_output_port_net;
  out_3 <= reinterpret2_output_port_net;
  out_4 <= reinterpret3_output_port_net;
  out_5 <= reinterpret4_output_port_net;
  out_6 <= reinterpret5_output_port_net;
  out_7 <= reinterpret6_output_port_net;
  out_8 <= reinterpret7_output_port_net;
  out_9 <= reinterpret8_output_port_net;
  out_10 <= reinterpret9_output_port_net;
  out_11 <= reinterpret10_output_port_net;
  out_12 <= reinterpret11_output_port_net;
  out_13 <= reinterpret12_output_port_net;
  out_14 <= reinterpret13_output_port_net;
  out_15 <= reinterpret14_output_port_net;
  out_16 <= reinterpret15_output_port_net;
  slice0_y_net <= in_1;
  slice1_y_net <= in_2;
  slice2_y_net <= in_3;
  slice3_y_net <= in_4;
  slice4_y_net <= in_5;
  slice5_y_net <= in_6;
  slice6_y_net <= in_7;
  slice7_y_net <= in_8;
  slice8_y_net <= in_9;
  slice9_y_net <= in_10;
  slice10_y_net <= in_11;
  slice11_y_net <= in_12;
  slice12_y_net <= in_13;
  slice13_y_net <= in_14;
  slice14_y_net <= in_15;
  slice15_y_net <= in_16;
  reinterpret0 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice0_y_net,
    output_port => reinterpret0_output_port_net
  );
  reinterpret1 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice1_y_net,
    output_port => reinterpret1_output_port_net
  );
  reinterpret2 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice2_y_net,
    output_port => reinterpret2_output_port_net
  );
  reinterpret3 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice3_y_net,
    output_port => reinterpret3_output_port_net
  );
  reinterpret4 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice4_y_net,
    output_port => reinterpret4_output_port_net
  );
  reinterpret5 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice5_y_net,
    output_port => reinterpret5_output_port_net
  );
  reinterpret6 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice6_y_net,
    output_port => reinterpret6_output_port_net
  );
  reinterpret7 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice7_y_net,
    output_port => reinterpret7_output_port_net
  );
  reinterpret8 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice8_y_net,
    output_port => reinterpret8_output_port_net
  );
  reinterpret9 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice9_y_net,
    output_port => reinterpret9_output_port_net
  );
  reinterpret10 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice10_y_net,
    output_port => reinterpret10_output_port_net
  );
  reinterpret11 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice11_y_net,
    output_port => reinterpret11_output_port_net
  );
  reinterpret12 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice12_y_net,
    output_port => reinterpret12_output_port_net
  );
  reinterpret13 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice13_y_net,
    output_port => reinterpret13_output_port_net
  );
  reinterpret14 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice14_y_net,
    output_port => reinterpret14_output_port_net
  );
  reinterpret15 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice15_y_net,
    output_port => reinterpret15_output_port_net
  );
end structural;
-- Generated from Simulink block PSB3_0/reordering extending buffer imag_1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_reordering_extending_buffer_imag_1 is
  port (
    in_reset : in std_logic_vector( 1-1 downto 0 );
    input1 : in std_logic_vector( 16-1 downto 0 );
    input2 : in std_logic_vector( 16-1 downto 0 );
    in_tvalid : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    vec_output_1 : out std_logic_vector( 16-1 downto 0 );
    vec_output_2 : out std_logic_vector( 16-1 downto 0 );
    vec_output_3 : out std_logic_vector( 16-1 downto 0 );
    vec_output_4 : out std_logic_vector( 16-1 downto 0 );
    vec_output_5 : out std_logic_vector( 16-1 downto 0 );
    vec_output_6 : out std_logic_vector( 16-1 downto 0 );
    vec_output_7 : out std_logic_vector( 16-1 downto 0 );
    vec_output_8 : out std_logic_vector( 16-1 downto 0 );
    vec_output_9 : out std_logic_vector( 16-1 downto 0 );
    vec_output_10 : out std_logic_vector( 16-1 downto 0 );
    vec_output_11 : out std_logic_vector( 16-1 downto 0 );
    vec_output_12 : out std_logic_vector( 16-1 downto 0 );
    vec_output_13 : out std_logic_vector( 16-1 downto 0 );
    vec_output_14 : out std_logic_vector( 16-1 downto 0 );
    vec_output_15 : out std_logic_vector( 16-1 downto 0 );
    vec_output_16 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_reordering_extending_buffer_imag_1;
architecture structural of psb3_0_reordering_extending_buffer_imag_1 is 
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal gin_tl_reset_net : std_logic_vector( 1-1 downto 0 );
  signal mux0_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 16-1 downto 0 );
  signal delay19_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 16-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 1-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 16-1 downto 0 );
  signal ce_net : std_logic;
  signal slice4_y_net : std_logic_vector( 16-1 downto 0 );
  signal dual_port_ram_0_douta_net : std_logic_vector( 16-1 downto 0 );
  signal bitbasher_out_x0_net : std_logic_vector( 256-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 16-1 downto 0 );
  signal dual_port_ram_1_doutb_net : std_logic_vector( 16-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 16-1 downto 0 );
  signal dual_port_ram_0_doutb_net : std_logic_vector( 16-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 16-1 downto 0 );
  signal mux5_y_net : std_logic_vector( 256-1 downto 0 );
  signal dual_port_ram_1_douta_net : std_logic_vector( 16-1 downto 0 );
  signal constant_op_net : std_logic_vector( 1-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 16-1 downto 0 );
  signal clk_net : std_logic;
  signal constant2_op_net : std_logic_vector( 1-1 downto 0 );
  signal mux4_y_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal bitbasher1_out_x0_net : std_logic_vector( 256-1 downto 0 );
  signal single_port_ram_data_out_net : std_logic_vector( 1-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 9-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 9-1 downto 0 );
  signal odd_addr_w_op_net : std_logic_vector( 9-1 downto 0 );
  signal we_0 : std_logic_vector( 1-1 downto 0 );
  signal delay10_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay11_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 16-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 16-1 downto 0 );
  signal inverter_op_net : std_logic_vector( 1-1 downto 0 );
  signal even_addr_w_op_net : std_logic_vector( 9-1 downto 0 );
  signal mux2_y_net : std_logic_vector( 9-1 downto 0 );
  signal mux3_y_net : std_logic_vector( 9-1 downto 0 );
  signal delay9_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux4_y_net : std_logic_vector( 9-1 downto 0 );
  signal delay7_q_net : std_logic_vector( 8-1 downto 0 );
  signal addr_r_op_net : std_logic_vector( 8-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 9-1 downto 0 );
  signal addr_control_op_net : std_logic_vector( 9-1 downto 0 );
  signal out_in_1024_out_x0_net : std_logic_vector( 9-1 downto 0 );
begin
  vec_output_1 <= reinterpret0_output_port_net;
  vec_output_2 <= reinterpret1_output_port_net;
  vec_output_3 <= reinterpret2_output_port_net;
  vec_output_4 <= reinterpret3_output_port_net;
  vec_output_5 <= reinterpret4_output_port_net;
  vec_output_6 <= reinterpret5_output_port_net;
  vec_output_7 <= reinterpret6_output_port_net;
  vec_output_8 <= reinterpret7_output_port_net;
  vec_output_9 <= reinterpret8_output_port_net;
  vec_output_10 <= reinterpret9_output_port_net;
  vec_output_11 <= reinterpret10_output_port_net;
  vec_output_12 <= reinterpret11_output_port_net;
  vec_output_13 <= reinterpret12_output_port_net;
  vec_output_14 <= reinterpret13_output_port_net;
  vec_output_15 <= reinterpret14_output_port_net;
  vec_output_16 <= reinterpret15_output_port_net;
  gin_tl_reset_net <= in_reset;
  mux0_y_net <= input1;
  mux4_y_net_x0 <= input2;
  delay19_q_net <= in_tvalid;
  clk_net <= clk_1;
  ce_net <= ce_1;
  scalar_to_vector4 : entity xil_defaultlib.psb3_0_scalar_to_vector4_x0 
  port map (
    i => mux5_y_net,
    o_1 => slice0_y_net,
    o_2 => slice1_y_net,
    o_3 => slice2_y_net,
    o_4 => slice3_y_net,
    o_5 => slice4_y_net,
    o_6 => slice5_y_net,
    o_7 => slice6_y_net,
    o_8 => slice7_y_net,
    o_9 => slice8_y_net,
    o_10 => slice9_y_net,
    o_11 => slice10_y_net,
    o_12 => slice11_y_net,
    o_13 => slice12_y_net,
    o_14 => slice13_y_net,
    o_15 => slice14_y_net,
    o_16 => slice15_y_net
  );
  vector_reinterpret : entity xil_defaultlib.psb3_0_vector_reinterpret_x3 
  port map (
    in_1 => slice0_y_net,
    in_2 => slice1_y_net,
    in_3 => slice2_y_net,
    in_4 => slice3_y_net,
    in_5 => slice4_y_net,
    in_6 => slice5_y_net,
    in_7 => slice6_y_net,
    in_8 => slice7_y_net,
    in_9 => slice8_y_net,
    in_10 => slice9_y_net,
    in_11 => slice10_y_net,
    in_12 => slice11_y_net,
    in_13 => slice12_y_net,
    in_14 => slice13_y_net,
    in_15 => slice14_y_net,
    in_16 => slice15_y_net,
    out_1 => reinterpret0_output_port_net,
    out_2 => reinterpret1_output_port_net,
    out_3 => reinterpret2_output_port_net,
    out_4 => reinterpret3_output_port_net,
    out_5 => reinterpret4_output_port_net,
    out_6 => reinterpret5_output_port_net,
    out_7 => reinterpret6_output_port_net,
    out_8 => reinterpret7_output_port_net,
    out_9 => reinterpret8_output_port_net,
    out_10 => reinterpret9_output_port_net,
    out_11 => reinterpret10_output_port_net,
    out_12 => reinterpret11_output_port_net,
    out_13 => reinterpret12_output_port_net,
    out_14 => reinterpret13_output_port_net,
    out_15 => reinterpret14_output_port_net,
    out_16 => reinterpret15_output_port_net
  );
  bitbasher : entity xil_defaultlib.sysgen_bitbasher_4648460ba6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    a => dual_port_ram_0_douta_net,
    b => dual_port_ram_0_doutb_net,
    out_x0 => bitbasher_out_x0_net
  );
  bitbasher1 : entity xil_defaultlib.sysgen_bitbasher_4648460ba6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    a => dual_port_ram_1_douta_net,
    b => dual_port_ram_1_doutb_net,
    out_x0 => bitbasher1_out_x0_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_de9059c03f 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_71e89d757c 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  constant2 : entity xil_defaultlib.sysgen_constant_71e89d757c 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant2_op_net
  );
  delay : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => single_port_ram_data_out_net,
    clk => clk_net,
    ce => ce_net,
    q => we_0
  );
  delay1 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 16
  )
  port map (
    en => '1',
    rst => '0',
    d => mux0_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay10 : entity xil_defaultlib.sysgen_delay_906db00812 
  port map (
    clr => '0',
    d => constant1_op_net,
    rst => gin_tl_reset_net,
    clk => clk_net,
    ce => ce_net,
    q => delay10_q_net
  );
  delay11 : entity xil_defaultlib.sysgen_delay_906db00812 
  port map (
    clr => '0',
    d => constant2_op_net,
    rst => gin_tl_reset_net,
    clk => clk_net,
    ce => ce_net,
    q => delay11_q_net
  );
  delay2 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 16
  )
  port map (
    en => '1',
    rst => '0',
    d => mux4_y_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay3 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => we_0,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  delay4 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => inverter_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net
  );
  delay5 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 9
  )
  port map (
    en => '1',
    rst => '0',
    d => even_addr_w_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  delay6 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 9
  )
  port map (
    en => '1',
    rst => '0',
    d => odd_addr_w_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay6_q_net
  );
  delay7 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 8
  )
  port map (
    en => '1',
    rst => '0',
    d => addr_r_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay7_q_net
  );
  delay9 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay9_q_net
  );
  dual_port_ram_0 : entity xil_defaultlib.psb3_0_xltdpram 
  generic map (
    addr_width_b => 9,
    clocking_mode => "common_clock",
    data_width_b => 16,
    latency => 1,
    mem_init_file => "xpm_c5fd30_vivado.mem",
    mem_size => 8192,
    mem_type => "block",
    read_reset_a => "0",
    read_reset_b => "0",
    width => 16,
    width_addr => 9,
    write_mode_a => "read_first",
    write_mode_b => "read_first"
  )
  port map (
    ena => "1",
    rsta => "0",
    rstb => "0",
    addra => mux1_y_net,
    dina => delay1_q_net,
    wea => delay3_q_net,
    addrb => mux2_y_net,
    dinb => delay2_q_net,
    web => delay3_q_net,
    enb => delay11_q_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dual_port_ram_0_douta_net,
    doutb => dual_port_ram_0_doutb_net
  );
  dual_port_ram_1 : entity xil_defaultlib.psb3_0_xltdpram 
  generic map (
    addr_width_b => 9,
    clocking_mode => "common_clock",
    data_width_b => 16,
    latency => 1,
    mem_init_file => "xpm_c5fd30_vivado.mem",
    mem_size => 8192,
    mem_type => "block",
    read_reset_a => "0",
    read_reset_b => "0",
    width => 16,
    width_addr => 9,
    write_mode_a => "read_first",
    write_mode_b => "read_first"
  )
  port map (
    ena => "1",
    rsta => "0",
    rstb => "0",
    addra => mux3_y_net,
    dina => delay1_q_net,
    wea => delay4_q_net,
    addrb => mux4_y_net,
    dinb => delay2_q_net,
    web => delay4_q_net,
    enb => delay10_q_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dual_port_ram_1_douta_net,
    doutb => dual_port_ram_1_doutb_net
  );
  inverter : entity xil_defaultlib.sysgen_inverter_ac5174c184 
  port map (
    clr => '0',
    ip => single_port_ram_data_out_net,
    clk => clk_net,
    ce => ce_net,
    op => inverter_op_net
  );
  mux1 : entity xil_defaultlib.sysgen_mux_303302b1e4 
  port map (
    clr => '0',
    sel => we_0,
    d0 => delay7_q_net,
    d1 => delay5_q_net,
    clk => clk_net,
    ce => ce_net,
    y => mux1_y_net
  );
  mux2 : entity xil_defaultlib.sysgen_mux_c7d0cfa098 
  port map (
    clr => '0',
    sel => we_0,
    d0 => out_in_1024_out_x0_net,
    d1 => delay6_q_net,
    clk => clk_net,
    ce => ce_net,
    y => mux2_y_net
  );
  mux3 : entity xil_defaultlib.sysgen_mux_303302b1e4 
  port map (
    clr => '0',
    sel => inverter_op_net,
    d0 => delay7_q_net,
    d1 => delay5_q_net,
    clk => clk_net,
    ce => ce_net,
    y => mux3_y_net
  );
  mux4 : entity xil_defaultlib.sysgen_mux_c7d0cfa098 
  port map (
    clr => '0',
    sel => inverter_op_net,
    d0 => out_in_1024_out_x0_net,
    d1 => delay6_q_net,
    clk => clk_net,
    ce => ce_net,
    y => mux4_y_net
  );
  mux5 : entity xil_defaultlib.sysgen_mux_1f606cf16b 
  port map (
    clr => '0',
    sel => delay9_q_net,
    d0 => bitbasher_out_x0_net,
    d1 => bitbasher1_out_x0_net,
    clk => clk_net,
    ce => ce_net,
    y => mux5_y_net
  );
  single_port_ram : entity xil_defaultlib.psb3_0_xlspram 
  generic map (
    init_value => b"0",
    latency => 1,
    mem_init_file => "xpm_95b604_vivado.mem",
    mem_size => 512,
    mem_type => "block",
    read_reset_val => "0",
    width => 1,
    width_addr => 9,
    write_mode_a => "read_first",
    xpm_lat => 1
  )
  port map (
    en => "1",
    rst => "0",
    addr => addr_control_op_net,
    data_in => constant_op_net,
    we => constant_op_net,
    clk => clk_net,
    ce => ce_net,
    data_out => single_port_ram_data_out_net
  );
  addr_control : entity xil_defaultlib.psb3_0_xlcounter_free 
  generic map (
    core_name0 => "psb3_0_c_counter_binary_v12_0_i4",
    op_arith => xlUnsigned,
    op_width => 9
  )
  port map (
    clr => '0',
    rst => gin_tl_reset_net,
    en => delay19_q_net,
    clk => clk_net,
    ce => ce_net,
    op => addr_control_op_net
  );
  addr_r : entity xil_defaultlib.psb3_0_xlcounter_free 
  generic map (
    core_name0 => "psb3_0_c_counter_binary_v12_0_i3",
    op_arith => xlUnsigned,
    op_width => 8
  )
  port map (
    clr => '0',
    rst => gin_tl_reset_net,
    en => delay19_q_net,
    clk => clk_net,
    ce => ce_net,
    op => addr_r_op_net
  );
  even_addr_w : entity xil_defaultlib.psb3_0_xlcounter_free 
  generic map (
    core_name0 => "psb3_0_c_counter_binary_v12_0_i5",
    op_arith => xlUnsigned,
    op_width => 9
  )
  port map (
    clr => '0',
    rst => gin_tl_reset_net,
    en => delay19_q_net,
    clk => clk_net,
    ce => ce_net,
    op => even_addr_w_op_net
  );
  odd_addr_w : entity xil_defaultlib.psb3_0_xlcounter_free 
  generic map (
    core_name0 => "psb3_0_c_counter_binary_v12_0_i6",
    op_arith => xlUnsigned,
    op_width => 9
  )
  port map (
    clr => '0',
    rst => gin_tl_reset_net,
    en => delay19_q_net,
    clk => clk_net,
    ce => ce_net,
    op => odd_addr_w_op_net
  );
  out_in_1024 : entity xil_defaultlib.sysgen_bitbasher_a62d2ce679 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in_x0 => delay7_q_net,
    out_x0 => out_in_1024_out_x0_net
  );
end structural;
-- Generated from Simulink block PSB3_0/reordering extending buffer imag_2/Scalar to Vector4
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_scalar_to_vector4_x1 is
  port (
    i : in std_logic_vector( 256-1 downto 0 );
    o_1 : out std_logic_vector( 16-1 downto 0 );
    o_2 : out std_logic_vector( 16-1 downto 0 );
    o_3 : out std_logic_vector( 16-1 downto 0 );
    o_4 : out std_logic_vector( 16-1 downto 0 );
    o_5 : out std_logic_vector( 16-1 downto 0 );
    o_6 : out std_logic_vector( 16-1 downto 0 );
    o_7 : out std_logic_vector( 16-1 downto 0 );
    o_8 : out std_logic_vector( 16-1 downto 0 );
    o_9 : out std_logic_vector( 16-1 downto 0 );
    o_10 : out std_logic_vector( 16-1 downto 0 );
    o_11 : out std_logic_vector( 16-1 downto 0 );
    o_12 : out std_logic_vector( 16-1 downto 0 );
    o_13 : out std_logic_vector( 16-1 downto 0 );
    o_14 : out std_logic_vector( 16-1 downto 0 );
    o_15 : out std_logic_vector( 16-1 downto 0 );
    o_16 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_scalar_to_vector4_x1;
architecture structural of psb3_0_scalar_to_vector4_x1 is 
  signal slice1_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 16-1 downto 0 );
  signal mux5_y_net : std_logic_vector( 256-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 16-1 downto 0 );
begin
  o_1 <= slice0_y_net;
  o_2 <= slice1_y_net;
  o_3 <= slice2_y_net;
  o_4 <= slice3_y_net;
  o_5 <= slice4_y_net;
  o_6 <= slice5_y_net;
  o_7 <= slice6_y_net;
  o_8 <= slice7_y_net;
  o_9 <= slice8_y_net;
  o_10 <= slice9_y_net;
  o_11 <= slice10_y_net;
  o_12 <= slice11_y_net;
  o_13 <= slice12_y_net;
  o_14 <= slice13_y_net;
  o_15 <= slice14_y_net;
  o_16 <= slice15_y_net;
  mux5_y_net <= i;
  slice0 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 15,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice0_y_net
  );
  slice1 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 16,
    new_msb => 31,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice1_y_net
  );
  slice2 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 32,
    new_msb => 47,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice2_y_net
  );
  slice3 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 48,
    new_msb => 63,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice3_y_net
  );
  slice4 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 64,
    new_msb => 79,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice4_y_net
  );
  slice5 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 80,
    new_msb => 95,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice5_y_net
  );
  slice6 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 96,
    new_msb => 111,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice6_y_net
  );
  slice7 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 112,
    new_msb => 127,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice7_y_net
  );
  slice8 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 128,
    new_msb => 143,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice8_y_net
  );
  slice9 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 144,
    new_msb => 159,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice9_y_net
  );
  slice10 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 160,
    new_msb => 175,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice10_y_net
  );
  slice11 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 176,
    new_msb => 191,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice11_y_net
  );
  slice12 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 192,
    new_msb => 207,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice12_y_net
  );
  slice13 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 208,
    new_msb => 223,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice13_y_net
  );
  slice14 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 224,
    new_msb => 239,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice14_y_net
  );
  slice15 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 240,
    new_msb => 255,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice15_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/reordering extending buffer imag_2/Vector Reinterpret
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_reinterpret_x4 is
  port (
    in_1 : in std_logic_vector( 16-1 downto 0 );
    in_2 : in std_logic_vector( 16-1 downto 0 );
    in_3 : in std_logic_vector( 16-1 downto 0 );
    in_4 : in std_logic_vector( 16-1 downto 0 );
    in_5 : in std_logic_vector( 16-1 downto 0 );
    in_6 : in std_logic_vector( 16-1 downto 0 );
    in_7 : in std_logic_vector( 16-1 downto 0 );
    in_8 : in std_logic_vector( 16-1 downto 0 );
    in_9 : in std_logic_vector( 16-1 downto 0 );
    in_10 : in std_logic_vector( 16-1 downto 0 );
    in_11 : in std_logic_vector( 16-1 downto 0 );
    in_12 : in std_logic_vector( 16-1 downto 0 );
    in_13 : in std_logic_vector( 16-1 downto 0 );
    in_14 : in std_logic_vector( 16-1 downto 0 );
    in_15 : in std_logic_vector( 16-1 downto 0 );
    in_16 : in std_logic_vector( 16-1 downto 0 );
    out_1 : out std_logic_vector( 16-1 downto 0 );
    out_2 : out std_logic_vector( 16-1 downto 0 );
    out_3 : out std_logic_vector( 16-1 downto 0 );
    out_4 : out std_logic_vector( 16-1 downto 0 );
    out_5 : out std_logic_vector( 16-1 downto 0 );
    out_6 : out std_logic_vector( 16-1 downto 0 );
    out_7 : out std_logic_vector( 16-1 downto 0 );
    out_8 : out std_logic_vector( 16-1 downto 0 );
    out_9 : out std_logic_vector( 16-1 downto 0 );
    out_10 : out std_logic_vector( 16-1 downto 0 );
    out_11 : out std_logic_vector( 16-1 downto 0 );
    out_12 : out std_logic_vector( 16-1 downto 0 );
    out_13 : out std_logic_vector( 16-1 downto 0 );
    out_14 : out std_logic_vector( 16-1 downto 0 );
    out_15 : out std_logic_vector( 16-1 downto 0 );
    out_16 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_vector_reinterpret_x4;
architecture structural of psb3_0_vector_reinterpret_x4 is 
  signal slice8_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 16-1 downto 0 );
begin
  out_1 <= reinterpret0_output_port_net;
  out_2 <= reinterpret1_output_port_net;
  out_3 <= reinterpret2_output_port_net;
  out_4 <= reinterpret3_output_port_net;
  out_5 <= reinterpret4_output_port_net;
  out_6 <= reinterpret5_output_port_net;
  out_7 <= reinterpret6_output_port_net;
  out_8 <= reinterpret7_output_port_net;
  out_9 <= reinterpret8_output_port_net;
  out_10 <= reinterpret9_output_port_net;
  out_11 <= reinterpret10_output_port_net;
  out_12 <= reinterpret11_output_port_net;
  out_13 <= reinterpret12_output_port_net;
  out_14 <= reinterpret13_output_port_net;
  out_15 <= reinterpret14_output_port_net;
  out_16 <= reinterpret15_output_port_net;
  slice0_y_net <= in_1;
  slice1_y_net <= in_2;
  slice2_y_net <= in_3;
  slice3_y_net <= in_4;
  slice4_y_net <= in_5;
  slice5_y_net <= in_6;
  slice6_y_net <= in_7;
  slice7_y_net <= in_8;
  slice8_y_net <= in_9;
  slice9_y_net <= in_10;
  slice10_y_net <= in_11;
  slice11_y_net <= in_12;
  slice12_y_net <= in_13;
  slice13_y_net <= in_14;
  slice14_y_net <= in_15;
  slice15_y_net <= in_16;
  reinterpret0 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice0_y_net,
    output_port => reinterpret0_output_port_net
  );
  reinterpret1 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice1_y_net,
    output_port => reinterpret1_output_port_net
  );
  reinterpret2 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice2_y_net,
    output_port => reinterpret2_output_port_net
  );
  reinterpret3 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice3_y_net,
    output_port => reinterpret3_output_port_net
  );
  reinterpret4 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice4_y_net,
    output_port => reinterpret4_output_port_net
  );
  reinterpret5 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice5_y_net,
    output_port => reinterpret5_output_port_net
  );
  reinterpret6 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice6_y_net,
    output_port => reinterpret6_output_port_net
  );
  reinterpret7 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice7_y_net,
    output_port => reinterpret7_output_port_net
  );
  reinterpret8 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice8_y_net,
    output_port => reinterpret8_output_port_net
  );
  reinterpret9 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice9_y_net,
    output_port => reinterpret9_output_port_net
  );
  reinterpret10 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice10_y_net,
    output_port => reinterpret10_output_port_net
  );
  reinterpret11 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice11_y_net,
    output_port => reinterpret11_output_port_net
  );
  reinterpret12 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice12_y_net,
    output_port => reinterpret12_output_port_net
  );
  reinterpret13 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice13_y_net,
    output_port => reinterpret13_output_port_net
  );
  reinterpret14 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice14_y_net,
    output_port => reinterpret14_output_port_net
  );
  reinterpret15 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice15_y_net,
    output_port => reinterpret15_output_port_net
  );
end structural;
-- Generated from Simulink block PSB3_0/reordering extending buffer imag_2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_reordering_extending_buffer_imag_2 is
  port (
    in_reset : in std_logic_vector( 1-1 downto 0 );
    input1 : in std_logic_vector( 16-1 downto 0 );
    input2 : in std_logic_vector( 16-1 downto 0 );
    in_tvalid : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    vec_output_1 : out std_logic_vector( 16-1 downto 0 );
    vec_output_2 : out std_logic_vector( 16-1 downto 0 );
    vec_output_3 : out std_logic_vector( 16-1 downto 0 );
    vec_output_4 : out std_logic_vector( 16-1 downto 0 );
    vec_output_5 : out std_logic_vector( 16-1 downto 0 );
    vec_output_6 : out std_logic_vector( 16-1 downto 0 );
    vec_output_7 : out std_logic_vector( 16-1 downto 0 );
    vec_output_8 : out std_logic_vector( 16-1 downto 0 );
    vec_output_9 : out std_logic_vector( 16-1 downto 0 );
    vec_output_10 : out std_logic_vector( 16-1 downto 0 );
    vec_output_11 : out std_logic_vector( 16-1 downto 0 );
    vec_output_12 : out std_logic_vector( 16-1 downto 0 );
    vec_output_13 : out std_logic_vector( 16-1 downto 0 );
    vec_output_14 : out std_logic_vector( 16-1 downto 0 );
    vec_output_15 : out std_logic_vector( 16-1 downto 0 );
    vec_output_16 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_reordering_extending_buffer_imag_2;
architecture structural of psb3_0_reordering_extending_buffer_imag_2 is 
  signal delay3_q_net : std_logic_vector( 1-1 downto 0 );
  signal inverter_op_net : std_logic_vector( 1-1 downto 0 );
  signal odd_addr_w_op_net : std_logic_vector( 9-1 downto 0 );
  signal delay7_q_net : std_logic_vector( 8-1 downto 0 );
  signal addr_r_op_net : std_logic_vector( 8-1 downto 0 );
  signal delay11_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 16-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 9-1 downto 0 );
  signal even_addr_w_op_net : std_logic_vector( 9-1 downto 0 );
  signal delay10_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 16-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 9-1 downto 0 );
  signal delay9_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux2_y_net : std_logic_vector( 9-1 downto 0 );
  signal mux3_y_net : std_logic_vector( 9-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 9-1 downto 0 );
  signal mux4_y_net : std_logic_vector( 9-1 downto 0 );
  signal out_in_1024_out_x0_net : std_logic_vector( 9-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mux5_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal gin_tl_reset_net : std_logic_vector( 1-1 downto 0 );
  signal delay19_q_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal mux1_y_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal ce_net : std_logic;
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 16-1 downto 0 );
  signal mux5_y_net_x0 : std_logic_vector( 256-1 downto 0 );
  signal we_0 : std_logic_vector( 1-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 16-1 downto 0 );
  signal bitbasher1_out_x0_net : std_logic_vector( 256-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 16-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 1-1 downto 0 );
  signal dual_port_ram_0_doutb_net : std_logic_vector( 16-1 downto 0 );
  signal constant2_op_net : std_logic_vector( 1-1 downto 0 );
  signal single_port_ram_data_out_net : std_logic_vector( 1-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 16-1 downto 0 );
  signal dual_port_ram_0_douta_net : std_logic_vector( 16-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 16-1 downto 0 );
  signal constant_op_net : std_logic_vector( 1-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 16-1 downto 0 );
  signal bitbasher_out_x0_net : std_logic_vector( 256-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 16-1 downto 0 );
  signal dual_port_ram_1_douta_net : std_logic_vector( 16-1 downto 0 );
  signal dual_port_ram_1_doutb_net : std_logic_vector( 16-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 16-1 downto 0 );
  signal addr_control_op_net : std_logic_vector( 9-1 downto 0 );
begin
  vec_output_1 <= reinterpret0_output_port_net;
  vec_output_2 <= reinterpret1_output_port_net;
  vec_output_3 <= reinterpret2_output_port_net;
  vec_output_4 <= reinterpret3_output_port_net;
  vec_output_5 <= reinterpret4_output_port_net;
  vec_output_6 <= reinterpret5_output_port_net;
  vec_output_7 <= reinterpret6_output_port_net;
  vec_output_8 <= reinterpret7_output_port_net;
  vec_output_9 <= reinterpret8_output_port_net;
  vec_output_10 <= reinterpret9_output_port_net;
  vec_output_11 <= reinterpret10_output_port_net;
  vec_output_12 <= reinterpret11_output_port_net;
  vec_output_13 <= reinterpret12_output_port_net;
  vec_output_14 <= reinterpret13_output_port_net;
  vec_output_15 <= reinterpret14_output_port_net;
  vec_output_16 <= reinterpret15_output_port_net;
  gin_tl_reset_net <= in_reset;
  mux1_y_net_x0 <= input1;
  mux5_y_net <= input2;
  delay19_q_net <= in_tvalid;
  clk_net <= clk_1;
  ce_net <= ce_1;
  scalar_to_vector4 : entity xil_defaultlib.psb3_0_scalar_to_vector4_x1 
  port map (
    i => mux5_y_net_x0,
    o_1 => slice0_y_net,
    o_2 => slice1_y_net,
    o_3 => slice2_y_net,
    o_4 => slice3_y_net,
    o_5 => slice4_y_net,
    o_6 => slice5_y_net,
    o_7 => slice6_y_net,
    o_8 => slice7_y_net,
    o_9 => slice8_y_net,
    o_10 => slice9_y_net,
    o_11 => slice10_y_net,
    o_12 => slice11_y_net,
    o_13 => slice12_y_net,
    o_14 => slice13_y_net,
    o_15 => slice14_y_net,
    o_16 => slice15_y_net
  );
  vector_reinterpret : entity xil_defaultlib.psb3_0_vector_reinterpret_x4 
  port map (
    in_1 => slice0_y_net,
    in_2 => slice1_y_net,
    in_3 => slice2_y_net,
    in_4 => slice3_y_net,
    in_5 => slice4_y_net,
    in_6 => slice5_y_net,
    in_7 => slice6_y_net,
    in_8 => slice7_y_net,
    in_9 => slice8_y_net,
    in_10 => slice9_y_net,
    in_11 => slice10_y_net,
    in_12 => slice11_y_net,
    in_13 => slice12_y_net,
    in_14 => slice13_y_net,
    in_15 => slice14_y_net,
    in_16 => slice15_y_net,
    out_1 => reinterpret0_output_port_net,
    out_2 => reinterpret1_output_port_net,
    out_3 => reinterpret2_output_port_net,
    out_4 => reinterpret3_output_port_net,
    out_5 => reinterpret4_output_port_net,
    out_6 => reinterpret5_output_port_net,
    out_7 => reinterpret6_output_port_net,
    out_8 => reinterpret7_output_port_net,
    out_9 => reinterpret8_output_port_net,
    out_10 => reinterpret9_output_port_net,
    out_11 => reinterpret10_output_port_net,
    out_12 => reinterpret11_output_port_net,
    out_13 => reinterpret12_output_port_net,
    out_14 => reinterpret13_output_port_net,
    out_15 => reinterpret14_output_port_net,
    out_16 => reinterpret15_output_port_net
  );
  bitbasher : entity xil_defaultlib.sysgen_bitbasher_4648460ba6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    a => dual_port_ram_0_douta_net,
    b => dual_port_ram_0_doutb_net,
    out_x0 => bitbasher_out_x0_net
  );
  bitbasher1 : entity xil_defaultlib.sysgen_bitbasher_4648460ba6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    a => dual_port_ram_1_douta_net,
    b => dual_port_ram_1_doutb_net,
    out_x0 => bitbasher1_out_x0_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_de9059c03f 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_71e89d757c 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  constant2 : entity xil_defaultlib.sysgen_constant_71e89d757c 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant2_op_net
  );
  delay : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => single_port_ram_data_out_net,
    clk => clk_net,
    ce => ce_net,
    q => we_0
  );
  delay1 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 16
  )
  port map (
    en => '1',
    rst => '0',
    d => mux1_y_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay10 : entity xil_defaultlib.sysgen_delay_906db00812 
  port map (
    clr => '0',
    d => constant1_op_net,
    rst => gin_tl_reset_net,
    clk => clk_net,
    ce => ce_net,
    q => delay10_q_net
  );
  delay11 : entity xil_defaultlib.sysgen_delay_906db00812 
  port map (
    clr => '0',
    d => constant2_op_net,
    rst => gin_tl_reset_net,
    clk => clk_net,
    ce => ce_net,
    q => delay11_q_net
  );
  delay2 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 16
  )
  port map (
    en => '1',
    rst => '0',
    d => mux5_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay3 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => we_0,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  delay4 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => inverter_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net
  );
  delay5 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 9
  )
  port map (
    en => '1',
    rst => '0',
    d => even_addr_w_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  delay6 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 9
  )
  port map (
    en => '1',
    rst => '0',
    d => odd_addr_w_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay6_q_net
  );
  delay7 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 8
  )
  port map (
    en => '1',
    rst => '0',
    d => addr_r_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay7_q_net
  );
  delay9 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay9_q_net
  );
  dual_port_ram_0 : entity xil_defaultlib.psb3_0_xltdpram 
  generic map (
    addr_width_b => 9,
    clocking_mode => "common_clock",
    data_width_b => 16,
    latency => 1,
    mem_init_file => "xpm_c5fd30_vivado.mem",
    mem_size => 8192,
    mem_type => "block",
    read_reset_a => "0",
    read_reset_b => "0",
    width => 16,
    width_addr => 9,
    write_mode_a => "read_first",
    write_mode_b => "read_first"
  )
  port map (
    ena => "1",
    rsta => "0",
    rstb => "0",
    addra => mux1_y_net,
    dina => delay1_q_net,
    wea => delay3_q_net,
    addrb => mux2_y_net,
    dinb => delay2_q_net,
    web => delay3_q_net,
    enb => delay11_q_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dual_port_ram_0_douta_net,
    doutb => dual_port_ram_0_doutb_net
  );
  dual_port_ram_1 : entity xil_defaultlib.psb3_0_xltdpram 
  generic map (
    addr_width_b => 9,
    clocking_mode => "common_clock",
    data_width_b => 16,
    latency => 1,
    mem_init_file => "xpm_c5fd30_vivado.mem",
    mem_size => 8192,
    mem_type => "block",
    read_reset_a => "0",
    read_reset_b => "0",
    width => 16,
    width_addr => 9,
    write_mode_a => "read_first",
    write_mode_b => "read_first"
  )
  port map (
    ena => "1",
    rsta => "0",
    rstb => "0",
    addra => mux3_y_net,
    dina => delay1_q_net,
    wea => delay4_q_net,
    addrb => mux4_y_net,
    dinb => delay2_q_net,
    web => delay4_q_net,
    enb => delay10_q_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dual_port_ram_1_douta_net,
    doutb => dual_port_ram_1_doutb_net
  );
  inverter : entity xil_defaultlib.sysgen_inverter_ac5174c184 
  port map (
    clr => '0',
    ip => single_port_ram_data_out_net,
    clk => clk_net,
    ce => ce_net,
    op => inverter_op_net
  );
  mux1 : entity xil_defaultlib.sysgen_mux_303302b1e4 
  port map (
    clr => '0',
    sel => we_0,
    d0 => delay7_q_net,
    d1 => delay5_q_net,
    clk => clk_net,
    ce => ce_net,
    y => mux1_y_net
  );
  mux2 : entity xil_defaultlib.sysgen_mux_c7d0cfa098 
  port map (
    clr => '0',
    sel => we_0,
    d0 => out_in_1024_out_x0_net,
    d1 => delay6_q_net,
    clk => clk_net,
    ce => ce_net,
    y => mux2_y_net
  );
  mux3 : entity xil_defaultlib.sysgen_mux_303302b1e4 
  port map (
    clr => '0',
    sel => inverter_op_net,
    d0 => delay7_q_net,
    d1 => delay5_q_net,
    clk => clk_net,
    ce => ce_net,
    y => mux3_y_net
  );
  mux4 : entity xil_defaultlib.sysgen_mux_c7d0cfa098 
  port map (
    clr => '0',
    sel => inverter_op_net,
    d0 => out_in_1024_out_x0_net,
    d1 => delay6_q_net,
    clk => clk_net,
    ce => ce_net,
    y => mux4_y_net
  );
  mux5 : entity xil_defaultlib.sysgen_mux_1f606cf16b 
  port map (
    clr => '0',
    sel => delay9_q_net,
    d0 => bitbasher_out_x0_net,
    d1 => bitbasher1_out_x0_net,
    clk => clk_net,
    ce => ce_net,
    y => mux5_y_net_x0
  );
  single_port_ram : entity xil_defaultlib.psb3_0_xlspram 
  generic map (
    init_value => b"0",
    latency => 1,
    mem_init_file => "xpm_95b604_vivado.mem",
    mem_size => 512,
    mem_type => "block",
    read_reset_val => "0",
    width => 1,
    width_addr => 9,
    write_mode_a => "read_first",
    xpm_lat => 1
  )
  port map (
    en => "1",
    rst => "0",
    addr => addr_control_op_net,
    data_in => constant_op_net,
    we => constant_op_net,
    clk => clk_net,
    ce => ce_net,
    data_out => single_port_ram_data_out_net
  );
  addr_control : entity xil_defaultlib.psb3_0_xlcounter_free 
  generic map (
    core_name0 => "psb3_0_c_counter_binary_v12_0_i4",
    op_arith => xlUnsigned,
    op_width => 9
  )
  port map (
    clr => '0',
    rst => gin_tl_reset_net,
    en => delay19_q_net,
    clk => clk_net,
    ce => ce_net,
    op => addr_control_op_net
  );
  addr_r : entity xil_defaultlib.psb3_0_xlcounter_free 
  generic map (
    core_name0 => "psb3_0_c_counter_binary_v12_0_i3",
    op_arith => xlUnsigned,
    op_width => 8
  )
  port map (
    clr => '0',
    rst => gin_tl_reset_net,
    en => delay19_q_net,
    clk => clk_net,
    ce => ce_net,
    op => addr_r_op_net
  );
  even_addr_w : entity xil_defaultlib.psb3_0_xlcounter_free 
  generic map (
    core_name0 => "psb3_0_c_counter_binary_v12_0_i5",
    op_arith => xlUnsigned,
    op_width => 9
  )
  port map (
    clr => '0',
    rst => gin_tl_reset_net,
    en => delay19_q_net,
    clk => clk_net,
    ce => ce_net,
    op => even_addr_w_op_net
  );
  odd_addr_w : entity xil_defaultlib.psb3_0_xlcounter_free 
  generic map (
    core_name0 => "psb3_0_c_counter_binary_v12_0_i6",
    op_arith => xlUnsigned,
    op_width => 9
  )
  port map (
    clr => '0',
    rst => gin_tl_reset_net,
    en => delay19_q_net,
    clk => clk_net,
    ce => ce_net,
    op => odd_addr_w_op_net
  );
  out_in_1024 : entity xil_defaultlib.sysgen_bitbasher_a62d2ce679 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in_x0 => delay7_q_net,
    out_x0 => out_in_1024_out_x0_net
  );
end structural;
-- Generated from Simulink block PSB3_0/reordering extending buffer imag_3/Scalar to Vector4
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_scalar_to_vector4_x2 is
  port (
    i : in std_logic_vector( 256-1 downto 0 );
    o_1 : out std_logic_vector( 16-1 downto 0 );
    o_2 : out std_logic_vector( 16-1 downto 0 );
    o_3 : out std_logic_vector( 16-1 downto 0 );
    o_4 : out std_logic_vector( 16-1 downto 0 );
    o_5 : out std_logic_vector( 16-1 downto 0 );
    o_6 : out std_logic_vector( 16-1 downto 0 );
    o_7 : out std_logic_vector( 16-1 downto 0 );
    o_8 : out std_logic_vector( 16-1 downto 0 );
    o_9 : out std_logic_vector( 16-1 downto 0 );
    o_10 : out std_logic_vector( 16-1 downto 0 );
    o_11 : out std_logic_vector( 16-1 downto 0 );
    o_12 : out std_logic_vector( 16-1 downto 0 );
    o_13 : out std_logic_vector( 16-1 downto 0 );
    o_14 : out std_logic_vector( 16-1 downto 0 );
    o_15 : out std_logic_vector( 16-1 downto 0 );
    o_16 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_scalar_to_vector4_x2;
architecture structural of psb3_0_scalar_to_vector4_x2 is 
  signal slice0_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 16-1 downto 0 );
  signal mux5_y_net : std_logic_vector( 256-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 16-1 downto 0 );
begin
  o_1 <= slice0_y_net;
  o_2 <= slice1_y_net;
  o_3 <= slice2_y_net;
  o_4 <= slice3_y_net;
  o_5 <= slice4_y_net;
  o_6 <= slice5_y_net;
  o_7 <= slice6_y_net;
  o_8 <= slice7_y_net;
  o_9 <= slice8_y_net;
  o_10 <= slice9_y_net;
  o_11 <= slice10_y_net;
  o_12 <= slice11_y_net;
  o_13 <= slice12_y_net;
  o_14 <= slice13_y_net;
  o_15 <= slice14_y_net;
  o_16 <= slice15_y_net;
  mux5_y_net <= i;
  slice0 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 15,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice0_y_net
  );
  slice1 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 16,
    new_msb => 31,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice1_y_net
  );
  slice2 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 32,
    new_msb => 47,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice2_y_net
  );
  slice3 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 48,
    new_msb => 63,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice3_y_net
  );
  slice4 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 64,
    new_msb => 79,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice4_y_net
  );
  slice5 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 80,
    new_msb => 95,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice5_y_net
  );
  slice6 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 96,
    new_msb => 111,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice6_y_net
  );
  slice7 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 112,
    new_msb => 127,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice7_y_net
  );
  slice8 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 128,
    new_msb => 143,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice8_y_net
  );
  slice9 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 144,
    new_msb => 159,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice9_y_net
  );
  slice10 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 160,
    new_msb => 175,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice10_y_net
  );
  slice11 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 176,
    new_msb => 191,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice11_y_net
  );
  slice12 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 192,
    new_msb => 207,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice12_y_net
  );
  slice13 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 208,
    new_msb => 223,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice13_y_net
  );
  slice14 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 224,
    new_msb => 239,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice14_y_net
  );
  slice15 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 240,
    new_msb => 255,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice15_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/reordering extending buffer imag_3/Vector Reinterpret
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_reinterpret_x5 is
  port (
    in_1 : in std_logic_vector( 16-1 downto 0 );
    in_2 : in std_logic_vector( 16-1 downto 0 );
    in_3 : in std_logic_vector( 16-1 downto 0 );
    in_4 : in std_logic_vector( 16-1 downto 0 );
    in_5 : in std_logic_vector( 16-1 downto 0 );
    in_6 : in std_logic_vector( 16-1 downto 0 );
    in_7 : in std_logic_vector( 16-1 downto 0 );
    in_8 : in std_logic_vector( 16-1 downto 0 );
    in_9 : in std_logic_vector( 16-1 downto 0 );
    in_10 : in std_logic_vector( 16-1 downto 0 );
    in_11 : in std_logic_vector( 16-1 downto 0 );
    in_12 : in std_logic_vector( 16-1 downto 0 );
    in_13 : in std_logic_vector( 16-1 downto 0 );
    in_14 : in std_logic_vector( 16-1 downto 0 );
    in_15 : in std_logic_vector( 16-1 downto 0 );
    in_16 : in std_logic_vector( 16-1 downto 0 );
    out_1 : out std_logic_vector( 16-1 downto 0 );
    out_2 : out std_logic_vector( 16-1 downto 0 );
    out_3 : out std_logic_vector( 16-1 downto 0 );
    out_4 : out std_logic_vector( 16-1 downto 0 );
    out_5 : out std_logic_vector( 16-1 downto 0 );
    out_6 : out std_logic_vector( 16-1 downto 0 );
    out_7 : out std_logic_vector( 16-1 downto 0 );
    out_8 : out std_logic_vector( 16-1 downto 0 );
    out_9 : out std_logic_vector( 16-1 downto 0 );
    out_10 : out std_logic_vector( 16-1 downto 0 );
    out_11 : out std_logic_vector( 16-1 downto 0 );
    out_12 : out std_logic_vector( 16-1 downto 0 );
    out_13 : out std_logic_vector( 16-1 downto 0 );
    out_14 : out std_logic_vector( 16-1 downto 0 );
    out_15 : out std_logic_vector( 16-1 downto 0 );
    out_16 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_vector_reinterpret_x5;
architecture structural of psb3_0_vector_reinterpret_x5 is 
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 16-1 downto 0 );
begin
  out_1 <= reinterpret0_output_port_net;
  out_2 <= reinterpret1_output_port_net;
  out_3 <= reinterpret2_output_port_net;
  out_4 <= reinterpret3_output_port_net;
  out_5 <= reinterpret4_output_port_net;
  out_6 <= reinterpret5_output_port_net;
  out_7 <= reinterpret6_output_port_net;
  out_8 <= reinterpret7_output_port_net;
  out_9 <= reinterpret8_output_port_net;
  out_10 <= reinterpret9_output_port_net;
  out_11 <= reinterpret10_output_port_net;
  out_12 <= reinterpret11_output_port_net;
  out_13 <= reinterpret12_output_port_net;
  out_14 <= reinterpret13_output_port_net;
  out_15 <= reinterpret14_output_port_net;
  out_16 <= reinterpret15_output_port_net;
  slice0_y_net <= in_1;
  slice1_y_net <= in_2;
  slice2_y_net <= in_3;
  slice3_y_net <= in_4;
  slice4_y_net <= in_5;
  slice5_y_net <= in_6;
  slice6_y_net <= in_7;
  slice7_y_net <= in_8;
  slice8_y_net <= in_9;
  slice9_y_net <= in_10;
  slice10_y_net <= in_11;
  slice11_y_net <= in_12;
  slice12_y_net <= in_13;
  slice13_y_net <= in_14;
  slice14_y_net <= in_15;
  slice15_y_net <= in_16;
  reinterpret0 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice0_y_net,
    output_port => reinterpret0_output_port_net
  );
  reinterpret1 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice1_y_net,
    output_port => reinterpret1_output_port_net
  );
  reinterpret2 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice2_y_net,
    output_port => reinterpret2_output_port_net
  );
  reinterpret3 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice3_y_net,
    output_port => reinterpret3_output_port_net
  );
  reinterpret4 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice4_y_net,
    output_port => reinterpret4_output_port_net
  );
  reinterpret5 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice5_y_net,
    output_port => reinterpret5_output_port_net
  );
  reinterpret6 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice6_y_net,
    output_port => reinterpret6_output_port_net
  );
  reinterpret7 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice7_y_net,
    output_port => reinterpret7_output_port_net
  );
  reinterpret8 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice8_y_net,
    output_port => reinterpret8_output_port_net
  );
  reinterpret9 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice9_y_net,
    output_port => reinterpret9_output_port_net
  );
  reinterpret10 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice10_y_net,
    output_port => reinterpret10_output_port_net
  );
  reinterpret11 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice11_y_net,
    output_port => reinterpret11_output_port_net
  );
  reinterpret12 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice12_y_net,
    output_port => reinterpret12_output_port_net
  );
  reinterpret13 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice13_y_net,
    output_port => reinterpret13_output_port_net
  );
  reinterpret14 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice14_y_net,
    output_port => reinterpret14_output_port_net
  );
  reinterpret15 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice15_y_net,
    output_port => reinterpret15_output_port_net
  );
end structural;
-- Generated from Simulink block PSB3_0/reordering extending buffer imag_3
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_reordering_extending_buffer_imag_3 is
  port (
    in_reset : in std_logic_vector( 1-1 downto 0 );
    input1 : in std_logic_vector( 16-1 downto 0 );
    input2 : in std_logic_vector( 16-1 downto 0 );
    in_tvalid : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    vec_output_1 : out std_logic_vector( 16-1 downto 0 );
    vec_output_2 : out std_logic_vector( 16-1 downto 0 );
    vec_output_3 : out std_logic_vector( 16-1 downto 0 );
    vec_output_4 : out std_logic_vector( 16-1 downto 0 );
    vec_output_5 : out std_logic_vector( 16-1 downto 0 );
    vec_output_6 : out std_logic_vector( 16-1 downto 0 );
    vec_output_7 : out std_logic_vector( 16-1 downto 0 );
    vec_output_8 : out std_logic_vector( 16-1 downto 0 );
    vec_output_9 : out std_logic_vector( 16-1 downto 0 );
    vec_output_10 : out std_logic_vector( 16-1 downto 0 );
    vec_output_11 : out std_logic_vector( 16-1 downto 0 );
    vec_output_12 : out std_logic_vector( 16-1 downto 0 );
    vec_output_13 : out std_logic_vector( 16-1 downto 0 );
    vec_output_14 : out std_logic_vector( 16-1 downto 0 );
    vec_output_15 : out std_logic_vector( 16-1 downto 0 );
    vec_output_16 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_reordering_extending_buffer_imag_3;
architecture structural of psb3_0_reordering_extending_buffer_imag_3 is 
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal delay19_q_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal clk_net : std_logic;
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal gin_tl_reset_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal ce_net : std_logic;
  signal slice0_y_net : std_logic_vector( 16-1 downto 0 );
  signal mux6_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mux2_y_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 16-1 downto 0 );
  signal we_0 : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 16-1 downto 0 );
  signal mux5_y_net : std_logic_vector( 256-1 downto 0 );
  signal bitbasher_out_x0_net : std_logic_vector( 256-1 downto 0 );
  signal dual_port_ram_0_doutb_net : std_logic_vector( 16-1 downto 0 );
  signal bitbasher1_out_x0_net : std_logic_vector( 256-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 16-1 downto 0 );
  signal dual_port_ram_1_douta_net : std_logic_vector( 16-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 16-1 downto 0 );
  signal dual_port_ram_0_douta_net : std_logic_vector( 16-1 downto 0 );
  signal constant_op_net : std_logic_vector( 1-1 downto 0 );
  signal constant2_op_net : std_logic_vector( 1-1 downto 0 );
  signal dual_port_ram_1_doutb_net : std_logic_vector( 16-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 16-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 1-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 16-1 downto 0 );
  signal single_port_ram_data_out_net : std_logic_vector( 1-1 downto 0 );
  signal delay9_q_net : std_logic_vector( 1-1 downto 0 );
  signal even_addr_w_op_net : std_logic_vector( 9-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 16-1 downto 0 );
  signal odd_addr_w_op_net : std_logic_vector( 9-1 downto 0 );
  signal addr_r_op_net : std_logic_vector( 8-1 downto 0 );
  signal delay11_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 1-1 downto 0 );
  signal inverter_op_net : std_logic_vector( 1-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 9-1 downto 0 );
  signal delay7_q_net : std_logic_vector( 8-1 downto 0 );
  signal delay10_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 9-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 9-1 downto 0 );
  signal mux4_y_net : std_logic_vector( 9-1 downto 0 );
  signal mux2_y_net : std_logic_vector( 9-1 downto 0 );
  signal out_in_1024_out_x0_net : std_logic_vector( 9-1 downto 0 );
  signal mux3_y_net : std_logic_vector( 9-1 downto 0 );
  signal addr_control_op_net : std_logic_vector( 9-1 downto 0 );
begin
  vec_output_1 <= reinterpret0_output_port_net;
  vec_output_2 <= reinterpret1_output_port_net;
  vec_output_3 <= reinterpret2_output_port_net;
  vec_output_4 <= reinterpret3_output_port_net;
  vec_output_5 <= reinterpret4_output_port_net;
  vec_output_6 <= reinterpret5_output_port_net;
  vec_output_7 <= reinterpret6_output_port_net;
  vec_output_8 <= reinterpret7_output_port_net;
  vec_output_9 <= reinterpret8_output_port_net;
  vec_output_10 <= reinterpret9_output_port_net;
  vec_output_11 <= reinterpret10_output_port_net;
  vec_output_12 <= reinterpret11_output_port_net;
  vec_output_13 <= reinterpret12_output_port_net;
  vec_output_14 <= reinterpret13_output_port_net;
  vec_output_15 <= reinterpret14_output_port_net;
  vec_output_16 <= reinterpret15_output_port_net;
  gin_tl_reset_net <= in_reset;
  mux2_y_net_x0 <= input1;
  mux6_y_net <= input2;
  delay19_q_net <= in_tvalid;
  clk_net <= clk_1;
  ce_net <= ce_1;
  scalar_to_vector4 : entity xil_defaultlib.psb3_0_scalar_to_vector4_x2 
  port map (
    i => mux5_y_net,
    o_1 => slice0_y_net,
    o_2 => slice1_y_net,
    o_3 => slice2_y_net,
    o_4 => slice3_y_net,
    o_5 => slice4_y_net,
    o_6 => slice5_y_net,
    o_7 => slice6_y_net,
    o_8 => slice7_y_net,
    o_9 => slice8_y_net,
    o_10 => slice9_y_net,
    o_11 => slice10_y_net,
    o_12 => slice11_y_net,
    o_13 => slice12_y_net,
    o_14 => slice13_y_net,
    o_15 => slice14_y_net,
    o_16 => slice15_y_net
  );
  vector_reinterpret : entity xil_defaultlib.psb3_0_vector_reinterpret_x5 
  port map (
    in_1 => slice0_y_net,
    in_2 => slice1_y_net,
    in_3 => slice2_y_net,
    in_4 => slice3_y_net,
    in_5 => slice4_y_net,
    in_6 => slice5_y_net,
    in_7 => slice6_y_net,
    in_8 => slice7_y_net,
    in_9 => slice8_y_net,
    in_10 => slice9_y_net,
    in_11 => slice10_y_net,
    in_12 => slice11_y_net,
    in_13 => slice12_y_net,
    in_14 => slice13_y_net,
    in_15 => slice14_y_net,
    in_16 => slice15_y_net,
    out_1 => reinterpret0_output_port_net,
    out_2 => reinterpret1_output_port_net,
    out_3 => reinterpret2_output_port_net,
    out_4 => reinterpret3_output_port_net,
    out_5 => reinterpret4_output_port_net,
    out_6 => reinterpret5_output_port_net,
    out_7 => reinterpret6_output_port_net,
    out_8 => reinterpret7_output_port_net,
    out_9 => reinterpret8_output_port_net,
    out_10 => reinterpret9_output_port_net,
    out_11 => reinterpret10_output_port_net,
    out_12 => reinterpret11_output_port_net,
    out_13 => reinterpret12_output_port_net,
    out_14 => reinterpret13_output_port_net,
    out_15 => reinterpret14_output_port_net,
    out_16 => reinterpret15_output_port_net
  );
  bitbasher : entity xil_defaultlib.sysgen_bitbasher_4648460ba6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    a => dual_port_ram_0_douta_net,
    b => dual_port_ram_0_doutb_net,
    out_x0 => bitbasher_out_x0_net
  );
  bitbasher1 : entity xil_defaultlib.sysgen_bitbasher_4648460ba6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    a => dual_port_ram_1_douta_net,
    b => dual_port_ram_1_doutb_net,
    out_x0 => bitbasher1_out_x0_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_de9059c03f 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_71e89d757c 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  constant2 : entity xil_defaultlib.sysgen_constant_71e89d757c 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant2_op_net
  );
  delay : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => single_port_ram_data_out_net,
    clk => clk_net,
    ce => ce_net,
    q => we_0
  );
  delay1 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 16
  )
  port map (
    en => '1',
    rst => '0',
    d => mux2_y_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay10 : entity xil_defaultlib.sysgen_delay_906db00812 
  port map (
    clr => '0',
    d => constant1_op_net,
    rst => gin_tl_reset_net,
    clk => clk_net,
    ce => ce_net,
    q => delay10_q_net
  );
  delay11 : entity xil_defaultlib.sysgen_delay_906db00812 
  port map (
    clr => '0',
    d => constant2_op_net,
    rst => gin_tl_reset_net,
    clk => clk_net,
    ce => ce_net,
    q => delay11_q_net
  );
  delay2 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 16
  )
  port map (
    en => '1',
    rst => '0',
    d => mux6_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay3 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => we_0,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  delay4 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => inverter_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net
  );
  delay5 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 9
  )
  port map (
    en => '1',
    rst => '0',
    d => even_addr_w_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  delay6 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 9
  )
  port map (
    en => '1',
    rst => '0',
    d => odd_addr_w_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay6_q_net
  );
  delay7 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 8
  )
  port map (
    en => '1',
    rst => '0',
    d => addr_r_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay7_q_net
  );
  delay9 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay9_q_net
  );
  dual_port_ram_0 : entity xil_defaultlib.psb3_0_xltdpram 
  generic map (
    addr_width_b => 9,
    clocking_mode => "common_clock",
    data_width_b => 16,
    latency => 1,
    mem_init_file => "xpm_c5fd30_vivado.mem",
    mem_size => 8192,
    mem_type => "block",
    read_reset_a => "0",
    read_reset_b => "0",
    width => 16,
    width_addr => 9,
    write_mode_a => "read_first",
    write_mode_b => "read_first"
  )
  port map (
    ena => "1",
    rsta => "0",
    rstb => "0",
    addra => mux1_y_net,
    dina => delay1_q_net,
    wea => delay3_q_net,
    addrb => mux2_y_net,
    dinb => delay2_q_net,
    web => delay3_q_net,
    enb => delay11_q_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dual_port_ram_0_douta_net,
    doutb => dual_port_ram_0_doutb_net
  );
  dual_port_ram_1 : entity xil_defaultlib.psb3_0_xltdpram 
  generic map (
    addr_width_b => 9,
    clocking_mode => "common_clock",
    data_width_b => 16,
    latency => 1,
    mem_init_file => "xpm_c5fd30_vivado.mem",
    mem_size => 8192,
    mem_type => "block",
    read_reset_a => "0",
    read_reset_b => "0",
    width => 16,
    width_addr => 9,
    write_mode_a => "read_first",
    write_mode_b => "read_first"
  )
  port map (
    ena => "1",
    rsta => "0",
    rstb => "0",
    addra => mux3_y_net,
    dina => delay1_q_net,
    wea => delay4_q_net,
    addrb => mux4_y_net,
    dinb => delay2_q_net,
    web => delay4_q_net,
    enb => delay10_q_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dual_port_ram_1_douta_net,
    doutb => dual_port_ram_1_doutb_net
  );
  inverter : entity xil_defaultlib.sysgen_inverter_ac5174c184 
  port map (
    clr => '0',
    ip => single_port_ram_data_out_net,
    clk => clk_net,
    ce => ce_net,
    op => inverter_op_net
  );
  mux1 : entity xil_defaultlib.sysgen_mux_303302b1e4 
  port map (
    clr => '0',
    sel => we_0,
    d0 => delay7_q_net,
    d1 => delay5_q_net,
    clk => clk_net,
    ce => ce_net,
    y => mux1_y_net
  );
  mux2 : entity xil_defaultlib.sysgen_mux_c7d0cfa098 
  port map (
    clr => '0',
    sel => we_0,
    d0 => out_in_1024_out_x0_net,
    d1 => delay6_q_net,
    clk => clk_net,
    ce => ce_net,
    y => mux2_y_net
  );
  mux3 : entity xil_defaultlib.sysgen_mux_303302b1e4 
  port map (
    clr => '0',
    sel => inverter_op_net,
    d0 => delay7_q_net,
    d1 => delay5_q_net,
    clk => clk_net,
    ce => ce_net,
    y => mux3_y_net
  );
  mux4 : entity xil_defaultlib.sysgen_mux_c7d0cfa098 
  port map (
    clr => '0',
    sel => inverter_op_net,
    d0 => out_in_1024_out_x0_net,
    d1 => delay6_q_net,
    clk => clk_net,
    ce => ce_net,
    y => mux4_y_net
  );
  mux5 : entity xil_defaultlib.sysgen_mux_1f606cf16b 
  port map (
    clr => '0',
    sel => delay9_q_net,
    d0 => bitbasher_out_x0_net,
    d1 => bitbasher1_out_x0_net,
    clk => clk_net,
    ce => ce_net,
    y => mux5_y_net
  );
  single_port_ram : entity xil_defaultlib.psb3_0_xlspram 
  generic map (
    init_value => b"0",
    latency => 1,
    mem_init_file => "xpm_95b604_vivado.mem",
    mem_size => 512,
    mem_type => "block",
    read_reset_val => "0",
    width => 1,
    width_addr => 9,
    write_mode_a => "read_first",
    xpm_lat => 1
  )
  port map (
    en => "1",
    rst => "0",
    addr => addr_control_op_net,
    data_in => constant_op_net,
    we => constant_op_net,
    clk => clk_net,
    ce => ce_net,
    data_out => single_port_ram_data_out_net
  );
  addr_control : entity xil_defaultlib.psb3_0_xlcounter_free 
  generic map (
    core_name0 => "psb3_0_c_counter_binary_v12_0_i4",
    op_arith => xlUnsigned,
    op_width => 9
  )
  port map (
    clr => '0',
    rst => gin_tl_reset_net,
    en => delay19_q_net,
    clk => clk_net,
    ce => ce_net,
    op => addr_control_op_net
  );
  addr_r : entity xil_defaultlib.psb3_0_xlcounter_free 
  generic map (
    core_name0 => "psb3_0_c_counter_binary_v12_0_i3",
    op_arith => xlUnsigned,
    op_width => 8
  )
  port map (
    clr => '0',
    rst => gin_tl_reset_net,
    en => delay19_q_net,
    clk => clk_net,
    ce => ce_net,
    op => addr_r_op_net
  );
  even_addr_w : entity xil_defaultlib.psb3_0_xlcounter_free 
  generic map (
    core_name0 => "psb3_0_c_counter_binary_v12_0_i5",
    op_arith => xlUnsigned,
    op_width => 9
  )
  port map (
    clr => '0',
    rst => gin_tl_reset_net,
    en => delay19_q_net,
    clk => clk_net,
    ce => ce_net,
    op => even_addr_w_op_net
  );
  odd_addr_w : entity xil_defaultlib.psb3_0_xlcounter_free 
  generic map (
    core_name0 => "psb3_0_c_counter_binary_v12_0_i6",
    op_arith => xlUnsigned,
    op_width => 9
  )
  port map (
    clr => '0',
    rst => gin_tl_reset_net,
    en => delay19_q_net,
    clk => clk_net,
    ce => ce_net,
    op => odd_addr_w_op_net
  );
  out_in_1024 : entity xil_defaultlib.sysgen_bitbasher_a62d2ce679 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in_x0 => delay7_q_net,
    out_x0 => out_in_1024_out_x0_net
  );
end structural;
-- Generated from Simulink block PSB3_0/reordering extending buffer imag_4/Scalar to Vector4
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_scalar_to_vector4_x3 is
  port (
    i : in std_logic_vector( 256-1 downto 0 );
    o_1 : out std_logic_vector( 16-1 downto 0 );
    o_2 : out std_logic_vector( 16-1 downto 0 );
    o_3 : out std_logic_vector( 16-1 downto 0 );
    o_4 : out std_logic_vector( 16-1 downto 0 );
    o_5 : out std_logic_vector( 16-1 downto 0 );
    o_6 : out std_logic_vector( 16-1 downto 0 );
    o_7 : out std_logic_vector( 16-1 downto 0 );
    o_8 : out std_logic_vector( 16-1 downto 0 );
    o_9 : out std_logic_vector( 16-1 downto 0 );
    o_10 : out std_logic_vector( 16-1 downto 0 );
    o_11 : out std_logic_vector( 16-1 downto 0 );
    o_12 : out std_logic_vector( 16-1 downto 0 );
    o_13 : out std_logic_vector( 16-1 downto 0 );
    o_14 : out std_logic_vector( 16-1 downto 0 );
    o_15 : out std_logic_vector( 16-1 downto 0 );
    o_16 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_scalar_to_vector4_x3;
architecture structural of psb3_0_scalar_to_vector4_x3 is 
  signal slice4_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 16-1 downto 0 );
  signal mux5_y_net : std_logic_vector( 256-1 downto 0 );
begin
  o_1 <= slice0_y_net;
  o_2 <= slice1_y_net;
  o_3 <= slice2_y_net;
  o_4 <= slice3_y_net;
  o_5 <= slice4_y_net;
  o_6 <= slice5_y_net;
  o_7 <= slice6_y_net;
  o_8 <= slice7_y_net;
  o_9 <= slice8_y_net;
  o_10 <= slice9_y_net;
  o_11 <= slice10_y_net;
  o_12 <= slice11_y_net;
  o_13 <= slice12_y_net;
  o_14 <= slice13_y_net;
  o_15 <= slice14_y_net;
  o_16 <= slice15_y_net;
  mux5_y_net <= i;
  slice0 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 15,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice0_y_net
  );
  slice1 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 16,
    new_msb => 31,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice1_y_net
  );
  slice2 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 32,
    new_msb => 47,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice2_y_net
  );
  slice3 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 48,
    new_msb => 63,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice3_y_net
  );
  slice4 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 64,
    new_msb => 79,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice4_y_net
  );
  slice5 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 80,
    new_msb => 95,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice5_y_net
  );
  slice6 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 96,
    new_msb => 111,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice6_y_net
  );
  slice7 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 112,
    new_msb => 127,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice7_y_net
  );
  slice8 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 128,
    new_msb => 143,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice8_y_net
  );
  slice9 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 144,
    new_msb => 159,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice9_y_net
  );
  slice10 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 160,
    new_msb => 175,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice10_y_net
  );
  slice11 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 176,
    new_msb => 191,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice11_y_net
  );
  slice12 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 192,
    new_msb => 207,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice12_y_net
  );
  slice13 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 208,
    new_msb => 223,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice13_y_net
  );
  slice14 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 224,
    new_msb => 239,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice14_y_net
  );
  slice15 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 240,
    new_msb => 255,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice15_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/reordering extending buffer imag_4/Vector Reinterpret
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_reinterpret_x6 is
  port (
    in_1 : in std_logic_vector( 16-1 downto 0 );
    in_2 : in std_logic_vector( 16-1 downto 0 );
    in_3 : in std_logic_vector( 16-1 downto 0 );
    in_4 : in std_logic_vector( 16-1 downto 0 );
    in_5 : in std_logic_vector( 16-1 downto 0 );
    in_6 : in std_logic_vector( 16-1 downto 0 );
    in_7 : in std_logic_vector( 16-1 downto 0 );
    in_8 : in std_logic_vector( 16-1 downto 0 );
    in_9 : in std_logic_vector( 16-1 downto 0 );
    in_10 : in std_logic_vector( 16-1 downto 0 );
    in_11 : in std_logic_vector( 16-1 downto 0 );
    in_12 : in std_logic_vector( 16-1 downto 0 );
    in_13 : in std_logic_vector( 16-1 downto 0 );
    in_14 : in std_logic_vector( 16-1 downto 0 );
    in_15 : in std_logic_vector( 16-1 downto 0 );
    in_16 : in std_logic_vector( 16-1 downto 0 );
    out_1 : out std_logic_vector( 16-1 downto 0 );
    out_2 : out std_logic_vector( 16-1 downto 0 );
    out_3 : out std_logic_vector( 16-1 downto 0 );
    out_4 : out std_logic_vector( 16-1 downto 0 );
    out_5 : out std_logic_vector( 16-1 downto 0 );
    out_6 : out std_logic_vector( 16-1 downto 0 );
    out_7 : out std_logic_vector( 16-1 downto 0 );
    out_8 : out std_logic_vector( 16-1 downto 0 );
    out_9 : out std_logic_vector( 16-1 downto 0 );
    out_10 : out std_logic_vector( 16-1 downto 0 );
    out_11 : out std_logic_vector( 16-1 downto 0 );
    out_12 : out std_logic_vector( 16-1 downto 0 );
    out_13 : out std_logic_vector( 16-1 downto 0 );
    out_14 : out std_logic_vector( 16-1 downto 0 );
    out_15 : out std_logic_vector( 16-1 downto 0 );
    out_16 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_vector_reinterpret_x6;
architecture structural of psb3_0_vector_reinterpret_x6 is 
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 16-1 downto 0 );
begin
  out_1 <= reinterpret0_output_port_net;
  out_2 <= reinterpret1_output_port_net;
  out_3 <= reinterpret2_output_port_net;
  out_4 <= reinterpret3_output_port_net;
  out_5 <= reinterpret4_output_port_net;
  out_6 <= reinterpret5_output_port_net;
  out_7 <= reinterpret6_output_port_net;
  out_8 <= reinterpret7_output_port_net;
  out_9 <= reinterpret8_output_port_net;
  out_10 <= reinterpret9_output_port_net;
  out_11 <= reinterpret10_output_port_net;
  out_12 <= reinterpret11_output_port_net;
  out_13 <= reinterpret12_output_port_net;
  out_14 <= reinterpret13_output_port_net;
  out_15 <= reinterpret14_output_port_net;
  out_16 <= reinterpret15_output_port_net;
  slice0_y_net <= in_1;
  slice1_y_net <= in_2;
  slice2_y_net <= in_3;
  slice3_y_net <= in_4;
  slice4_y_net <= in_5;
  slice5_y_net <= in_6;
  slice6_y_net <= in_7;
  slice7_y_net <= in_8;
  slice8_y_net <= in_9;
  slice9_y_net <= in_10;
  slice10_y_net <= in_11;
  slice11_y_net <= in_12;
  slice12_y_net <= in_13;
  slice13_y_net <= in_14;
  slice14_y_net <= in_15;
  slice15_y_net <= in_16;
  reinterpret0 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice0_y_net,
    output_port => reinterpret0_output_port_net
  );
  reinterpret1 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice1_y_net,
    output_port => reinterpret1_output_port_net
  );
  reinterpret2 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice2_y_net,
    output_port => reinterpret2_output_port_net
  );
  reinterpret3 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice3_y_net,
    output_port => reinterpret3_output_port_net
  );
  reinterpret4 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice4_y_net,
    output_port => reinterpret4_output_port_net
  );
  reinterpret5 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice5_y_net,
    output_port => reinterpret5_output_port_net
  );
  reinterpret6 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice6_y_net,
    output_port => reinterpret6_output_port_net
  );
  reinterpret7 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice7_y_net,
    output_port => reinterpret7_output_port_net
  );
  reinterpret8 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice8_y_net,
    output_port => reinterpret8_output_port_net
  );
  reinterpret9 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice9_y_net,
    output_port => reinterpret9_output_port_net
  );
  reinterpret10 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice10_y_net,
    output_port => reinterpret10_output_port_net
  );
  reinterpret11 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice11_y_net,
    output_port => reinterpret11_output_port_net
  );
  reinterpret12 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice12_y_net,
    output_port => reinterpret12_output_port_net
  );
  reinterpret13 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice13_y_net,
    output_port => reinterpret13_output_port_net
  );
  reinterpret14 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice14_y_net,
    output_port => reinterpret14_output_port_net
  );
  reinterpret15 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice15_y_net,
    output_port => reinterpret15_output_port_net
  );
end structural;
-- Generated from Simulink block PSB3_0/reordering extending buffer imag_4
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_reordering_extending_buffer_imag_4 is
  port (
    in_reset : in std_logic_vector( 1-1 downto 0 );
    input1 : in std_logic_vector( 16-1 downto 0 );
    input2 : in std_logic_vector( 16-1 downto 0 );
    in_tvalid : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    vec_output_1 : out std_logic_vector( 16-1 downto 0 );
    vec_output_2 : out std_logic_vector( 16-1 downto 0 );
    vec_output_3 : out std_logic_vector( 16-1 downto 0 );
    vec_output_4 : out std_logic_vector( 16-1 downto 0 );
    vec_output_5 : out std_logic_vector( 16-1 downto 0 );
    vec_output_6 : out std_logic_vector( 16-1 downto 0 );
    vec_output_7 : out std_logic_vector( 16-1 downto 0 );
    vec_output_8 : out std_logic_vector( 16-1 downto 0 );
    vec_output_9 : out std_logic_vector( 16-1 downto 0 );
    vec_output_10 : out std_logic_vector( 16-1 downto 0 );
    vec_output_11 : out std_logic_vector( 16-1 downto 0 );
    vec_output_12 : out std_logic_vector( 16-1 downto 0 );
    vec_output_13 : out std_logic_vector( 16-1 downto 0 );
    vec_output_14 : out std_logic_vector( 16-1 downto 0 );
    vec_output_15 : out std_logic_vector( 16-1 downto 0 );
    vec_output_16 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_reordering_extending_buffer_imag_4;
architecture structural of psb3_0_reordering_extending_buffer_imag_4 is 
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mux7_y_net : std_logic_vector( 16-1 downto 0 );
  signal clk_net : std_logic;
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 16-1 downto 0 );
  signal mux3_y_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 16-1 downto 0 );
  signal ce_net : std_logic;
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal gin_tl_reset_net : std_logic_vector( 1-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal delay19_q_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 16-1 downto 0 );
  signal constant2_op_net : std_logic_vector( 1-1 downto 0 );
  signal delay10_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 16-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 1-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 16-1 downto 0 );
  signal bitbasher1_out_x0_net : std_logic_vector( 256-1 downto 0 );
  signal dual_port_ram_1_doutb_net : std_logic_vector( 16-1 downto 0 );
  signal we_0 : std_logic_vector( 1-1 downto 0 );
  signal single_port_ram_data_out_net : std_logic_vector( 1-1 downto 0 );
  signal constant_op_net : std_logic_vector( 1-1 downto 0 );
  signal bitbasher_out_x0_net : std_logic_vector( 256-1 downto 0 );
  signal dual_port_ram_0_doutb_net : std_logic_vector( 16-1 downto 0 );
  signal dual_port_ram_0_douta_net : std_logic_vector( 16-1 downto 0 );
  signal dual_port_ram_1_douta_net : std_logic_vector( 16-1 downto 0 );
  signal mux5_y_net : std_logic_vector( 256-1 downto 0 );
  signal inverter_op_net : std_logic_vector( 1-1 downto 0 );
  signal even_addr_w_op_net : std_logic_vector( 9-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 16-1 downto 0 );
  signal addr_r_op_net : std_logic_vector( 8-1 downto 0 );
  signal delay11_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay9_q_net : std_logic_vector( 1-1 downto 0 );
  signal odd_addr_w_op_net : std_logic_vector( 9-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 9-1 downto 0 );
  signal delay7_q_net : std_logic_vector( 8-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 9-1 downto 0 );
  signal mux4_y_net : std_logic_vector( 9-1 downto 0 );
  signal mux2_y_net : std_logic_vector( 9-1 downto 0 );
  signal out_in_1024_out_x0_net : std_logic_vector( 9-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 9-1 downto 0 );
  signal mux3_y_net : std_logic_vector( 9-1 downto 0 );
  signal addr_control_op_net : std_logic_vector( 9-1 downto 0 );
begin
  vec_output_1 <= reinterpret0_output_port_net;
  vec_output_2 <= reinterpret1_output_port_net;
  vec_output_3 <= reinterpret2_output_port_net;
  vec_output_4 <= reinterpret3_output_port_net;
  vec_output_5 <= reinterpret4_output_port_net;
  vec_output_6 <= reinterpret5_output_port_net;
  vec_output_7 <= reinterpret6_output_port_net;
  vec_output_8 <= reinterpret7_output_port_net;
  vec_output_9 <= reinterpret8_output_port_net;
  vec_output_10 <= reinterpret9_output_port_net;
  vec_output_11 <= reinterpret10_output_port_net;
  vec_output_12 <= reinterpret11_output_port_net;
  vec_output_13 <= reinterpret12_output_port_net;
  vec_output_14 <= reinterpret13_output_port_net;
  vec_output_15 <= reinterpret14_output_port_net;
  vec_output_16 <= reinterpret15_output_port_net;
  gin_tl_reset_net <= in_reset;
  mux3_y_net_x0 <= input1;
  mux7_y_net <= input2;
  delay19_q_net <= in_tvalid;
  clk_net <= clk_1;
  ce_net <= ce_1;
  scalar_to_vector4 : entity xil_defaultlib.psb3_0_scalar_to_vector4_x3 
  port map (
    i => mux5_y_net,
    o_1 => slice0_y_net,
    o_2 => slice1_y_net,
    o_3 => slice2_y_net,
    o_4 => slice3_y_net,
    o_5 => slice4_y_net,
    o_6 => slice5_y_net,
    o_7 => slice6_y_net,
    o_8 => slice7_y_net,
    o_9 => slice8_y_net,
    o_10 => slice9_y_net,
    o_11 => slice10_y_net,
    o_12 => slice11_y_net,
    o_13 => slice12_y_net,
    o_14 => slice13_y_net,
    o_15 => slice14_y_net,
    o_16 => slice15_y_net
  );
  vector_reinterpret : entity xil_defaultlib.psb3_0_vector_reinterpret_x6 
  port map (
    in_1 => slice0_y_net,
    in_2 => slice1_y_net,
    in_3 => slice2_y_net,
    in_4 => slice3_y_net,
    in_5 => slice4_y_net,
    in_6 => slice5_y_net,
    in_7 => slice6_y_net,
    in_8 => slice7_y_net,
    in_9 => slice8_y_net,
    in_10 => slice9_y_net,
    in_11 => slice10_y_net,
    in_12 => slice11_y_net,
    in_13 => slice12_y_net,
    in_14 => slice13_y_net,
    in_15 => slice14_y_net,
    in_16 => slice15_y_net,
    out_1 => reinterpret0_output_port_net,
    out_2 => reinterpret1_output_port_net,
    out_3 => reinterpret2_output_port_net,
    out_4 => reinterpret3_output_port_net,
    out_5 => reinterpret4_output_port_net,
    out_6 => reinterpret5_output_port_net,
    out_7 => reinterpret6_output_port_net,
    out_8 => reinterpret7_output_port_net,
    out_9 => reinterpret8_output_port_net,
    out_10 => reinterpret9_output_port_net,
    out_11 => reinterpret10_output_port_net,
    out_12 => reinterpret11_output_port_net,
    out_13 => reinterpret12_output_port_net,
    out_14 => reinterpret13_output_port_net,
    out_15 => reinterpret14_output_port_net,
    out_16 => reinterpret15_output_port_net
  );
  bitbasher : entity xil_defaultlib.sysgen_bitbasher_4648460ba6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    a => dual_port_ram_0_douta_net,
    b => dual_port_ram_0_doutb_net,
    out_x0 => bitbasher_out_x0_net
  );
  bitbasher1 : entity xil_defaultlib.sysgen_bitbasher_4648460ba6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    a => dual_port_ram_1_douta_net,
    b => dual_port_ram_1_doutb_net,
    out_x0 => bitbasher1_out_x0_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_de9059c03f 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_71e89d757c 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  constant2 : entity xil_defaultlib.sysgen_constant_71e89d757c 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant2_op_net
  );
  delay : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => single_port_ram_data_out_net,
    clk => clk_net,
    ce => ce_net,
    q => we_0
  );
  delay1 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 16
  )
  port map (
    en => '1',
    rst => '0',
    d => mux3_y_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay10 : entity xil_defaultlib.sysgen_delay_906db00812 
  port map (
    clr => '0',
    d => constant1_op_net,
    rst => gin_tl_reset_net,
    clk => clk_net,
    ce => ce_net,
    q => delay10_q_net
  );
  delay11 : entity xil_defaultlib.sysgen_delay_906db00812 
  port map (
    clr => '0',
    d => constant2_op_net,
    rst => gin_tl_reset_net,
    clk => clk_net,
    ce => ce_net,
    q => delay11_q_net
  );
  delay2 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 16
  )
  port map (
    en => '1',
    rst => '0',
    d => mux7_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay3 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => we_0,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  delay4 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => inverter_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net
  );
  delay5 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 9
  )
  port map (
    en => '1',
    rst => '0',
    d => even_addr_w_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  delay6 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 9
  )
  port map (
    en => '1',
    rst => '0',
    d => odd_addr_w_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay6_q_net
  );
  delay7 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 8
  )
  port map (
    en => '1',
    rst => '0',
    d => addr_r_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay7_q_net
  );
  delay9 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay9_q_net
  );
  dual_port_ram_0 : entity xil_defaultlib.psb3_0_xltdpram 
  generic map (
    addr_width_b => 9,
    clocking_mode => "common_clock",
    data_width_b => 16,
    latency => 1,
    mem_init_file => "xpm_c5fd30_vivado.mem",
    mem_size => 8192,
    mem_type => "block",
    read_reset_a => "0",
    read_reset_b => "0",
    width => 16,
    width_addr => 9,
    write_mode_a => "read_first",
    write_mode_b => "read_first"
  )
  port map (
    ena => "1",
    rsta => "0",
    rstb => "0",
    addra => mux1_y_net,
    dina => delay1_q_net,
    wea => delay3_q_net,
    addrb => mux2_y_net,
    dinb => delay2_q_net,
    web => delay3_q_net,
    enb => delay11_q_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dual_port_ram_0_douta_net,
    doutb => dual_port_ram_0_doutb_net
  );
  dual_port_ram_1 : entity xil_defaultlib.psb3_0_xltdpram 
  generic map (
    addr_width_b => 9,
    clocking_mode => "common_clock",
    data_width_b => 16,
    latency => 1,
    mem_init_file => "xpm_c5fd30_vivado.mem",
    mem_size => 8192,
    mem_type => "block",
    read_reset_a => "0",
    read_reset_b => "0",
    width => 16,
    width_addr => 9,
    write_mode_a => "read_first",
    write_mode_b => "read_first"
  )
  port map (
    ena => "1",
    rsta => "0",
    rstb => "0",
    addra => mux3_y_net,
    dina => delay1_q_net,
    wea => delay4_q_net,
    addrb => mux4_y_net,
    dinb => delay2_q_net,
    web => delay4_q_net,
    enb => delay10_q_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dual_port_ram_1_douta_net,
    doutb => dual_port_ram_1_doutb_net
  );
  inverter : entity xil_defaultlib.sysgen_inverter_ac5174c184 
  port map (
    clr => '0',
    ip => single_port_ram_data_out_net,
    clk => clk_net,
    ce => ce_net,
    op => inverter_op_net
  );
  mux1 : entity xil_defaultlib.sysgen_mux_303302b1e4 
  port map (
    clr => '0',
    sel => we_0,
    d0 => delay7_q_net,
    d1 => delay5_q_net,
    clk => clk_net,
    ce => ce_net,
    y => mux1_y_net
  );
  mux2 : entity xil_defaultlib.sysgen_mux_c7d0cfa098 
  port map (
    clr => '0',
    sel => we_0,
    d0 => out_in_1024_out_x0_net,
    d1 => delay6_q_net,
    clk => clk_net,
    ce => ce_net,
    y => mux2_y_net
  );
  mux3 : entity xil_defaultlib.sysgen_mux_303302b1e4 
  port map (
    clr => '0',
    sel => inverter_op_net,
    d0 => delay7_q_net,
    d1 => delay5_q_net,
    clk => clk_net,
    ce => ce_net,
    y => mux3_y_net
  );
  mux4 : entity xil_defaultlib.sysgen_mux_c7d0cfa098 
  port map (
    clr => '0',
    sel => inverter_op_net,
    d0 => out_in_1024_out_x0_net,
    d1 => delay6_q_net,
    clk => clk_net,
    ce => ce_net,
    y => mux4_y_net
  );
  mux5 : entity xil_defaultlib.sysgen_mux_1f606cf16b 
  port map (
    clr => '0',
    sel => delay9_q_net,
    d0 => bitbasher_out_x0_net,
    d1 => bitbasher1_out_x0_net,
    clk => clk_net,
    ce => ce_net,
    y => mux5_y_net
  );
  single_port_ram : entity xil_defaultlib.psb3_0_xlspram 
  generic map (
    init_value => b"0",
    latency => 1,
    mem_init_file => "xpm_95b604_vivado.mem",
    mem_size => 512,
    mem_type => "block",
    read_reset_val => "0",
    width => 1,
    width_addr => 9,
    write_mode_a => "read_first",
    xpm_lat => 1
  )
  port map (
    en => "1",
    rst => "0",
    addr => addr_control_op_net,
    data_in => constant_op_net,
    we => constant_op_net,
    clk => clk_net,
    ce => ce_net,
    data_out => single_port_ram_data_out_net
  );
  addr_control : entity xil_defaultlib.psb3_0_xlcounter_free 
  generic map (
    core_name0 => "psb3_0_c_counter_binary_v12_0_i4",
    op_arith => xlUnsigned,
    op_width => 9
  )
  port map (
    clr => '0',
    rst => gin_tl_reset_net,
    en => delay19_q_net,
    clk => clk_net,
    ce => ce_net,
    op => addr_control_op_net
  );
  addr_r : entity xil_defaultlib.psb3_0_xlcounter_free 
  generic map (
    core_name0 => "psb3_0_c_counter_binary_v12_0_i3",
    op_arith => xlUnsigned,
    op_width => 8
  )
  port map (
    clr => '0',
    rst => gin_tl_reset_net,
    en => delay19_q_net,
    clk => clk_net,
    ce => ce_net,
    op => addr_r_op_net
  );
  even_addr_w : entity xil_defaultlib.psb3_0_xlcounter_free 
  generic map (
    core_name0 => "psb3_0_c_counter_binary_v12_0_i5",
    op_arith => xlUnsigned,
    op_width => 9
  )
  port map (
    clr => '0',
    rst => gin_tl_reset_net,
    en => delay19_q_net,
    clk => clk_net,
    ce => ce_net,
    op => even_addr_w_op_net
  );
  odd_addr_w : entity xil_defaultlib.psb3_0_xlcounter_free 
  generic map (
    core_name0 => "psb3_0_c_counter_binary_v12_0_i6",
    op_arith => xlUnsigned,
    op_width => 9
  )
  port map (
    clr => '0',
    rst => gin_tl_reset_net,
    en => delay19_q_net,
    clk => clk_net,
    ce => ce_net,
    op => odd_addr_w_op_net
  );
  out_in_1024 : entity xil_defaultlib.sysgen_bitbasher_a62d2ce679 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in_x0 => delay7_q_net,
    out_x0 => out_in_1024_out_x0_net
  );
end structural;
-- Generated from Simulink block PSB3_0/reordering extending buffer real_1/Scalar to Vector4
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_scalar_to_vector4_x4 is
  port (
    i : in std_logic_vector( 256-1 downto 0 );
    o_1 : out std_logic_vector( 16-1 downto 0 );
    o_2 : out std_logic_vector( 16-1 downto 0 );
    o_3 : out std_logic_vector( 16-1 downto 0 );
    o_4 : out std_logic_vector( 16-1 downto 0 );
    o_5 : out std_logic_vector( 16-1 downto 0 );
    o_6 : out std_logic_vector( 16-1 downto 0 );
    o_7 : out std_logic_vector( 16-1 downto 0 );
    o_8 : out std_logic_vector( 16-1 downto 0 );
    o_9 : out std_logic_vector( 16-1 downto 0 );
    o_10 : out std_logic_vector( 16-1 downto 0 );
    o_11 : out std_logic_vector( 16-1 downto 0 );
    o_12 : out std_logic_vector( 16-1 downto 0 );
    o_13 : out std_logic_vector( 16-1 downto 0 );
    o_14 : out std_logic_vector( 16-1 downto 0 );
    o_15 : out std_logic_vector( 16-1 downto 0 );
    o_16 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_scalar_to_vector4_x4;
architecture structural of psb3_0_scalar_to_vector4_x4 is 
  signal slice5_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 16-1 downto 0 );
  signal mux5_y_net : std_logic_vector( 256-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 16-1 downto 0 );
begin
  o_1 <= slice0_y_net;
  o_2 <= slice1_y_net;
  o_3 <= slice2_y_net;
  o_4 <= slice3_y_net;
  o_5 <= slice4_y_net;
  o_6 <= slice5_y_net;
  o_7 <= slice6_y_net;
  o_8 <= slice7_y_net;
  o_9 <= slice8_y_net;
  o_10 <= slice9_y_net;
  o_11 <= slice10_y_net;
  o_12 <= slice11_y_net;
  o_13 <= slice12_y_net;
  o_14 <= slice13_y_net;
  o_15 <= slice14_y_net;
  o_16 <= slice15_y_net;
  mux5_y_net <= i;
  slice0 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 15,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice0_y_net
  );
  slice1 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 16,
    new_msb => 31,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice1_y_net
  );
  slice2 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 32,
    new_msb => 47,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice2_y_net
  );
  slice3 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 48,
    new_msb => 63,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice3_y_net
  );
  slice4 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 64,
    new_msb => 79,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice4_y_net
  );
  slice5 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 80,
    new_msb => 95,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice5_y_net
  );
  slice6 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 96,
    new_msb => 111,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice6_y_net
  );
  slice7 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 112,
    new_msb => 127,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice7_y_net
  );
  slice8 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 128,
    new_msb => 143,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice8_y_net
  );
  slice9 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 144,
    new_msb => 159,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice9_y_net
  );
  slice10 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 160,
    new_msb => 175,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice10_y_net
  );
  slice11 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 176,
    new_msb => 191,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice11_y_net
  );
  slice12 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 192,
    new_msb => 207,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice12_y_net
  );
  slice13 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 208,
    new_msb => 223,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice13_y_net
  );
  slice14 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 224,
    new_msb => 239,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice14_y_net
  );
  slice15 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 240,
    new_msb => 255,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice15_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/reordering extending buffer real_1/Vector Reinterpret
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_reinterpret_x7 is
  port (
    in_1 : in std_logic_vector( 16-1 downto 0 );
    in_2 : in std_logic_vector( 16-1 downto 0 );
    in_3 : in std_logic_vector( 16-1 downto 0 );
    in_4 : in std_logic_vector( 16-1 downto 0 );
    in_5 : in std_logic_vector( 16-1 downto 0 );
    in_6 : in std_logic_vector( 16-1 downto 0 );
    in_7 : in std_logic_vector( 16-1 downto 0 );
    in_8 : in std_logic_vector( 16-1 downto 0 );
    in_9 : in std_logic_vector( 16-1 downto 0 );
    in_10 : in std_logic_vector( 16-1 downto 0 );
    in_11 : in std_logic_vector( 16-1 downto 0 );
    in_12 : in std_logic_vector( 16-1 downto 0 );
    in_13 : in std_logic_vector( 16-1 downto 0 );
    in_14 : in std_logic_vector( 16-1 downto 0 );
    in_15 : in std_logic_vector( 16-1 downto 0 );
    in_16 : in std_logic_vector( 16-1 downto 0 );
    out_1 : out std_logic_vector( 16-1 downto 0 );
    out_2 : out std_logic_vector( 16-1 downto 0 );
    out_3 : out std_logic_vector( 16-1 downto 0 );
    out_4 : out std_logic_vector( 16-1 downto 0 );
    out_5 : out std_logic_vector( 16-1 downto 0 );
    out_6 : out std_logic_vector( 16-1 downto 0 );
    out_7 : out std_logic_vector( 16-1 downto 0 );
    out_8 : out std_logic_vector( 16-1 downto 0 );
    out_9 : out std_logic_vector( 16-1 downto 0 );
    out_10 : out std_logic_vector( 16-1 downto 0 );
    out_11 : out std_logic_vector( 16-1 downto 0 );
    out_12 : out std_logic_vector( 16-1 downto 0 );
    out_13 : out std_logic_vector( 16-1 downto 0 );
    out_14 : out std_logic_vector( 16-1 downto 0 );
    out_15 : out std_logic_vector( 16-1 downto 0 );
    out_16 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_vector_reinterpret_x7;
architecture structural of psb3_0_vector_reinterpret_x7 is 
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 16-1 downto 0 );
begin
  out_1 <= reinterpret0_output_port_net;
  out_2 <= reinterpret1_output_port_net;
  out_3 <= reinterpret2_output_port_net;
  out_4 <= reinterpret3_output_port_net;
  out_5 <= reinterpret4_output_port_net;
  out_6 <= reinterpret5_output_port_net;
  out_7 <= reinterpret6_output_port_net;
  out_8 <= reinterpret7_output_port_net;
  out_9 <= reinterpret8_output_port_net;
  out_10 <= reinterpret9_output_port_net;
  out_11 <= reinterpret10_output_port_net;
  out_12 <= reinterpret11_output_port_net;
  out_13 <= reinterpret12_output_port_net;
  out_14 <= reinterpret13_output_port_net;
  out_15 <= reinterpret14_output_port_net;
  out_16 <= reinterpret15_output_port_net;
  slice0_y_net <= in_1;
  slice1_y_net <= in_2;
  slice2_y_net <= in_3;
  slice3_y_net <= in_4;
  slice4_y_net <= in_5;
  slice5_y_net <= in_6;
  slice6_y_net <= in_7;
  slice7_y_net <= in_8;
  slice8_y_net <= in_9;
  slice9_y_net <= in_10;
  slice10_y_net <= in_11;
  slice11_y_net <= in_12;
  slice12_y_net <= in_13;
  slice13_y_net <= in_14;
  slice14_y_net <= in_15;
  slice15_y_net <= in_16;
  reinterpret0 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice0_y_net,
    output_port => reinterpret0_output_port_net
  );
  reinterpret1 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice1_y_net,
    output_port => reinterpret1_output_port_net
  );
  reinterpret2 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice2_y_net,
    output_port => reinterpret2_output_port_net
  );
  reinterpret3 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice3_y_net,
    output_port => reinterpret3_output_port_net
  );
  reinterpret4 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice4_y_net,
    output_port => reinterpret4_output_port_net
  );
  reinterpret5 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice5_y_net,
    output_port => reinterpret5_output_port_net
  );
  reinterpret6 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice6_y_net,
    output_port => reinterpret6_output_port_net
  );
  reinterpret7 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice7_y_net,
    output_port => reinterpret7_output_port_net
  );
  reinterpret8 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice8_y_net,
    output_port => reinterpret8_output_port_net
  );
  reinterpret9 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice9_y_net,
    output_port => reinterpret9_output_port_net
  );
  reinterpret10 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice10_y_net,
    output_port => reinterpret10_output_port_net
  );
  reinterpret11 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice11_y_net,
    output_port => reinterpret11_output_port_net
  );
  reinterpret12 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice12_y_net,
    output_port => reinterpret12_output_port_net
  );
  reinterpret13 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice13_y_net,
    output_port => reinterpret13_output_port_net
  );
  reinterpret14 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice14_y_net,
    output_port => reinterpret14_output_port_net
  );
  reinterpret15 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice15_y_net,
    output_port => reinterpret15_output_port_net
  );
end structural;
-- Generated from Simulink block PSB3_0/reordering extending buffer real_1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_reordering_extending_buffer_real_1 is
  port (
    in_reset : in std_logic_vector( 1-1 downto 0 );
    input1 : in std_logic_vector( 16-1 downto 0 );
    input2 : in std_logic_vector( 16-1 downto 0 );
    in_tvalid : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    vec_output_1 : out std_logic_vector( 16-1 downto 0 );
    out_tvalid : out std_logic_vector( 1-1 downto 0 );
    vec_output_2 : out std_logic_vector( 16-1 downto 0 );
    vec_output_3 : out std_logic_vector( 16-1 downto 0 );
    vec_output_4 : out std_logic_vector( 16-1 downto 0 );
    vec_output_5 : out std_logic_vector( 16-1 downto 0 );
    vec_output_6 : out std_logic_vector( 16-1 downto 0 );
    vec_output_7 : out std_logic_vector( 16-1 downto 0 );
    vec_output_8 : out std_logic_vector( 16-1 downto 0 );
    vec_output_9 : out std_logic_vector( 16-1 downto 0 );
    vec_output_10 : out std_logic_vector( 16-1 downto 0 );
    vec_output_11 : out std_logic_vector( 16-1 downto 0 );
    vec_output_12 : out std_logic_vector( 16-1 downto 0 );
    vec_output_13 : out std_logic_vector( 16-1 downto 0 );
    vec_output_14 : out std_logic_vector( 16-1 downto 0 );
    vec_output_15 : out std_logic_vector( 16-1 downto 0 );
    vec_output_16 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_reordering_extending_buffer_real_1;
architecture structural of psb3_0_reordering_extending_buffer_real_1 is 
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal gin_tl_reset_net : std_logic_vector( 1-1 downto 0 );
  signal mux0_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal clk_net : std_logic;
  signal mux4_y_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal ce_net : std_logic;
  signal slice3_y_net : std_logic_vector( 16-1 downto 0 );
  signal delay19_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 16-1 downto 0 );
  signal mux5_y_net : std_logic_vector( 256-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 16-1 downto 0 );
  signal constant2_op_net : std_logic_vector( 1-1 downto 0 );
  signal we_0 : std_logic_vector( 1-1 downto 0 );
  signal bitbasher1_out_x0_net : std_logic_vector( 256-1 downto 0 );
  signal single_port_ram_data_out_net : std_logic_vector( 1-1 downto 0 );
  signal bitbasher_out_x0_net : std_logic_vector( 256-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 16-1 downto 0 );
  signal dual_port_ram_0_doutb_net : std_logic_vector( 16-1 downto 0 );
  signal constant_op_net : std_logic_vector( 1-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 1-1 downto 0 );
  signal dual_port_ram_1_doutb_net : std_logic_vector( 16-1 downto 0 );
  signal dual_port_ram_0_douta_net : std_logic_vector( 16-1 downto 0 );
  signal delay10_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay11_q_net : std_logic_vector( 1-1 downto 0 );
  signal dual_port_ram_1_douta_net : std_logic_vector( 16-1 downto 0 );
  signal odd_addr_w_op_net : std_logic_vector( 9-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 9-1 downto 0 );
  signal delay9_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay7_q_net : std_logic_vector( 8-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 16-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 9-1 downto 0 );
  signal inverter_op_net : std_logic_vector( 1-1 downto 0 );
  signal even_addr_w_op_net : std_logic_vector( 9-1 downto 0 );
  signal addr_r_op_net : std_logic_vector( 8-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux3_y_net : std_logic_vector( 9-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 9-1 downto 0 );
  signal mux2_y_net : std_logic_vector( 9-1 downto 0 );
  signal mux4_y_net : std_logic_vector( 9-1 downto 0 );
  signal out_in_1024_out_x0_net : std_logic_vector( 9-1 downto 0 );
  signal addr_control_op_net : std_logic_vector( 9-1 downto 0 );
begin
  vec_output_1 <= reinterpret0_output_port_net;
  out_tvalid <= delay8_q_net;
  vec_output_2 <= reinterpret1_output_port_net;
  vec_output_3 <= reinterpret2_output_port_net;
  vec_output_4 <= reinterpret3_output_port_net;
  vec_output_5 <= reinterpret4_output_port_net;
  vec_output_6 <= reinterpret5_output_port_net;
  vec_output_7 <= reinterpret6_output_port_net;
  vec_output_8 <= reinterpret7_output_port_net;
  vec_output_9 <= reinterpret8_output_port_net;
  vec_output_10 <= reinterpret9_output_port_net;
  vec_output_11 <= reinterpret10_output_port_net;
  vec_output_12 <= reinterpret11_output_port_net;
  vec_output_13 <= reinterpret12_output_port_net;
  vec_output_14 <= reinterpret13_output_port_net;
  vec_output_15 <= reinterpret14_output_port_net;
  vec_output_16 <= reinterpret15_output_port_net;
  gin_tl_reset_net <= in_reset;
  mux0_y_net <= input1;
  mux4_y_net_x0 <= input2;
  delay19_q_net <= in_tvalid;
  clk_net <= clk_1;
  ce_net <= ce_1;
  scalar_to_vector4 : entity xil_defaultlib.psb3_0_scalar_to_vector4_x4 
  port map (
    i => mux5_y_net,
    o_1 => slice0_y_net,
    o_2 => slice1_y_net,
    o_3 => slice2_y_net,
    o_4 => slice3_y_net,
    o_5 => slice4_y_net,
    o_6 => slice5_y_net,
    o_7 => slice6_y_net,
    o_8 => slice7_y_net,
    o_9 => slice8_y_net,
    o_10 => slice9_y_net,
    o_11 => slice10_y_net,
    o_12 => slice11_y_net,
    o_13 => slice12_y_net,
    o_14 => slice13_y_net,
    o_15 => slice14_y_net,
    o_16 => slice15_y_net
  );
  vector_reinterpret : entity xil_defaultlib.psb3_0_vector_reinterpret_x7 
  port map (
    in_1 => slice0_y_net,
    in_2 => slice1_y_net,
    in_3 => slice2_y_net,
    in_4 => slice3_y_net,
    in_5 => slice4_y_net,
    in_6 => slice5_y_net,
    in_7 => slice6_y_net,
    in_8 => slice7_y_net,
    in_9 => slice8_y_net,
    in_10 => slice9_y_net,
    in_11 => slice10_y_net,
    in_12 => slice11_y_net,
    in_13 => slice12_y_net,
    in_14 => slice13_y_net,
    in_15 => slice14_y_net,
    in_16 => slice15_y_net,
    out_1 => reinterpret0_output_port_net,
    out_2 => reinterpret1_output_port_net,
    out_3 => reinterpret2_output_port_net,
    out_4 => reinterpret3_output_port_net,
    out_5 => reinterpret4_output_port_net,
    out_6 => reinterpret5_output_port_net,
    out_7 => reinterpret6_output_port_net,
    out_8 => reinterpret7_output_port_net,
    out_9 => reinterpret8_output_port_net,
    out_10 => reinterpret9_output_port_net,
    out_11 => reinterpret10_output_port_net,
    out_12 => reinterpret11_output_port_net,
    out_13 => reinterpret12_output_port_net,
    out_14 => reinterpret13_output_port_net,
    out_15 => reinterpret14_output_port_net,
    out_16 => reinterpret15_output_port_net
  );
  bitbasher : entity xil_defaultlib.sysgen_bitbasher_4648460ba6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    a => dual_port_ram_0_douta_net,
    b => dual_port_ram_0_doutb_net,
    out_x0 => bitbasher_out_x0_net
  );
  bitbasher1 : entity xil_defaultlib.sysgen_bitbasher_4648460ba6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    a => dual_port_ram_1_douta_net,
    b => dual_port_ram_1_doutb_net,
    out_x0 => bitbasher1_out_x0_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_de9059c03f 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_71e89d757c 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  constant2 : entity xil_defaultlib.sysgen_constant_71e89d757c 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant2_op_net
  );
  delay : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => single_port_ram_data_out_net,
    clk => clk_net,
    ce => ce_net,
    q => we_0
  );
  delay1 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 16
  )
  port map (
    en => '1',
    rst => '0',
    d => mux0_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay10 : entity xil_defaultlib.sysgen_delay_906db00812 
  port map (
    clr => '0',
    d => constant1_op_net,
    rst => gin_tl_reset_net,
    clk => clk_net,
    ce => ce_net,
    q => delay10_q_net
  );
  delay11 : entity xil_defaultlib.sysgen_delay_906db00812 
  port map (
    clr => '0',
    d => constant2_op_net,
    rst => gin_tl_reset_net,
    clk => clk_net,
    ce => ce_net,
    q => delay11_q_net
  );
  delay2 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 16
  )
  port map (
    en => '1',
    rst => '0',
    d => mux4_y_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay3 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => we_0,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  delay4 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => inverter_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net
  );
  delay5 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 9
  )
  port map (
    en => '1',
    rst => '0',
    d => even_addr_w_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  delay6 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 9
  )
  port map (
    en => '1',
    rst => '0',
    d => odd_addr_w_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay6_q_net
  );
  delay7 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 8
  )
  port map (
    en => '1',
    rst => '0',
    d => addr_r_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay7_q_net
  );
  delay8 : entity xil_defaultlib.sysgen_delay_2c038b42f1 
  port map (
    clr => '0',
    d => delay19_q_net,
    rst => gin_tl_reset_net,
    clk => clk_net,
    ce => ce_net,
    q => delay8_q_net
  );
  delay9 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay9_q_net
  );
  dual_port_ram_0 : entity xil_defaultlib.psb3_0_xltdpram 
  generic map (
    addr_width_b => 9,
    clocking_mode => "common_clock",
    data_width_b => 16,
    latency => 1,
    mem_init_file => "xpm_c5fd30_vivado.mem",
    mem_size => 8192,
    mem_type => "block",
    read_reset_a => "0",
    read_reset_b => "0",
    width => 16,
    width_addr => 9,
    write_mode_a => "read_first",
    write_mode_b => "read_first"
  )
  port map (
    ena => "1",
    rsta => "0",
    rstb => "0",
    addra => mux1_y_net,
    dina => delay1_q_net,
    wea => delay3_q_net,
    addrb => mux2_y_net,
    dinb => delay2_q_net,
    web => delay3_q_net,
    enb => delay11_q_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dual_port_ram_0_douta_net,
    doutb => dual_port_ram_0_doutb_net
  );
  dual_port_ram_1 : entity xil_defaultlib.psb3_0_xltdpram 
  generic map (
    addr_width_b => 9,
    clocking_mode => "common_clock",
    data_width_b => 16,
    latency => 1,
    mem_init_file => "xpm_c5fd30_vivado.mem",
    mem_size => 8192,
    mem_type => "block",
    read_reset_a => "0",
    read_reset_b => "0",
    width => 16,
    width_addr => 9,
    write_mode_a => "read_first",
    write_mode_b => "read_first"
  )
  port map (
    ena => "1",
    rsta => "0",
    rstb => "0",
    addra => mux3_y_net,
    dina => delay1_q_net,
    wea => delay4_q_net,
    addrb => mux4_y_net,
    dinb => delay2_q_net,
    web => delay4_q_net,
    enb => delay10_q_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dual_port_ram_1_douta_net,
    doutb => dual_port_ram_1_doutb_net
  );
  inverter : entity xil_defaultlib.sysgen_inverter_ac5174c184 
  port map (
    clr => '0',
    ip => single_port_ram_data_out_net,
    clk => clk_net,
    ce => ce_net,
    op => inverter_op_net
  );
  mux1 : entity xil_defaultlib.sysgen_mux_303302b1e4 
  port map (
    clr => '0',
    sel => we_0,
    d0 => delay7_q_net,
    d1 => delay5_q_net,
    clk => clk_net,
    ce => ce_net,
    y => mux1_y_net
  );
  mux2 : entity xil_defaultlib.sysgen_mux_c7d0cfa098 
  port map (
    clr => '0',
    sel => we_0,
    d0 => out_in_1024_out_x0_net,
    d1 => delay6_q_net,
    clk => clk_net,
    ce => ce_net,
    y => mux2_y_net
  );
  mux3 : entity xil_defaultlib.sysgen_mux_303302b1e4 
  port map (
    clr => '0',
    sel => inverter_op_net,
    d0 => delay7_q_net,
    d1 => delay5_q_net,
    clk => clk_net,
    ce => ce_net,
    y => mux3_y_net
  );
  mux4 : entity xil_defaultlib.sysgen_mux_c7d0cfa098 
  port map (
    clr => '0',
    sel => inverter_op_net,
    d0 => out_in_1024_out_x0_net,
    d1 => delay6_q_net,
    clk => clk_net,
    ce => ce_net,
    y => mux4_y_net
  );
  mux5 : entity xil_defaultlib.sysgen_mux_1f606cf16b 
  port map (
    clr => '0',
    sel => delay9_q_net,
    d0 => bitbasher_out_x0_net,
    d1 => bitbasher1_out_x0_net,
    clk => clk_net,
    ce => ce_net,
    y => mux5_y_net
  );
  single_port_ram : entity xil_defaultlib.psb3_0_xlspram 
  generic map (
    init_value => b"0",
    latency => 1,
    mem_init_file => "xpm_95b604_vivado.mem",
    mem_size => 512,
    mem_type => "block",
    read_reset_val => "0",
    width => 1,
    width_addr => 9,
    write_mode_a => "read_first",
    xpm_lat => 1
  )
  port map (
    en => "1",
    rst => "0",
    addr => addr_control_op_net,
    data_in => constant_op_net,
    we => constant_op_net,
    clk => clk_net,
    ce => ce_net,
    data_out => single_port_ram_data_out_net
  );
  addr_control : entity xil_defaultlib.psb3_0_xlcounter_free 
  generic map (
    core_name0 => "psb3_0_c_counter_binary_v12_0_i4",
    op_arith => xlUnsigned,
    op_width => 9
  )
  port map (
    clr => '0',
    rst => gin_tl_reset_net,
    en => delay19_q_net,
    clk => clk_net,
    ce => ce_net,
    op => addr_control_op_net
  );
  addr_r : entity xil_defaultlib.psb3_0_xlcounter_free 
  generic map (
    core_name0 => "psb3_0_c_counter_binary_v12_0_i3",
    op_arith => xlUnsigned,
    op_width => 8
  )
  port map (
    clr => '0',
    rst => gin_tl_reset_net,
    en => delay19_q_net,
    clk => clk_net,
    ce => ce_net,
    op => addr_r_op_net
  );
  even_addr_w : entity xil_defaultlib.psb3_0_xlcounter_free 
  generic map (
    core_name0 => "psb3_0_c_counter_binary_v12_0_i5",
    op_arith => xlUnsigned,
    op_width => 9
  )
  port map (
    clr => '0',
    rst => gin_tl_reset_net,
    en => delay19_q_net,
    clk => clk_net,
    ce => ce_net,
    op => even_addr_w_op_net
  );
  odd_addr_w : entity xil_defaultlib.psb3_0_xlcounter_free 
  generic map (
    core_name0 => "psb3_0_c_counter_binary_v12_0_i6",
    op_arith => xlUnsigned,
    op_width => 9
  )
  port map (
    clr => '0',
    rst => gin_tl_reset_net,
    en => delay19_q_net,
    clk => clk_net,
    ce => ce_net,
    op => odd_addr_w_op_net
  );
  out_in_1024 : entity xil_defaultlib.sysgen_bitbasher_a62d2ce679 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in_x0 => delay7_q_net,
    out_x0 => out_in_1024_out_x0_net
  );
end structural;
-- Generated from Simulink block PSB3_0/reordering extending buffer real_2/Scalar to Vector4
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_scalar_to_vector4_x5 is
  port (
    i : in std_logic_vector( 256-1 downto 0 );
    o_1 : out std_logic_vector( 16-1 downto 0 );
    o_2 : out std_logic_vector( 16-1 downto 0 );
    o_3 : out std_logic_vector( 16-1 downto 0 );
    o_4 : out std_logic_vector( 16-1 downto 0 );
    o_5 : out std_logic_vector( 16-1 downto 0 );
    o_6 : out std_logic_vector( 16-1 downto 0 );
    o_7 : out std_logic_vector( 16-1 downto 0 );
    o_8 : out std_logic_vector( 16-1 downto 0 );
    o_9 : out std_logic_vector( 16-1 downto 0 );
    o_10 : out std_logic_vector( 16-1 downto 0 );
    o_11 : out std_logic_vector( 16-1 downto 0 );
    o_12 : out std_logic_vector( 16-1 downto 0 );
    o_13 : out std_logic_vector( 16-1 downto 0 );
    o_14 : out std_logic_vector( 16-1 downto 0 );
    o_15 : out std_logic_vector( 16-1 downto 0 );
    o_16 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_scalar_to_vector4_x5;
architecture structural of psb3_0_scalar_to_vector4_x5 is 
  signal slice4_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 16-1 downto 0 );
  signal mux5_y_net : std_logic_vector( 256-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 16-1 downto 0 );
begin
  o_1 <= slice0_y_net;
  o_2 <= slice1_y_net;
  o_3 <= slice2_y_net;
  o_4 <= slice3_y_net;
  o_5 <= slice4_y_net;
  o_6 <= slice5_y_net;
  o_7 <= slice6_y_net;
  o_8 <= slice7_y_net;
  o_9 <= slice8_y_net;
  o_10 <= slice9_y_net;
  o_11 <= slice10_y_net;
  o_12 <= slice11_y_net;
  o_13 <= slice12_y_net;
  o_14 <= slice13_y_net;
  o_15 <= slice14_y_net;
  o_16 <= slice15_y_net;
  mux5_y_net <= i;
  slice0 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 15,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice0_y_net
  );
  slice1 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 16,
    new_msb => 31,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice1_y_net
  );
  slice2 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 32,
    new_msb => 47,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice2_y_net
  );
  slice3 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 48,
    new_msb => 63,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice3_y_net
  );
  slice4 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 64,
    new_msb => 79,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice4_y_net
  );
  slice5 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 80,
    new_msb => 95,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice5_y_net
  );
  slice6 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 96,
    new_msb => 111,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice6_y_net
  );
  slice7 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 112,
    new_msb => 127,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice7_y_net
  );
  slice8 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 128,
    new_msb => 143,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice8_y_net
  );
  slice9 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 144,
    new_msb => 159,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice9_y_net
  );
  slice10 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 160,
    new_msb => 175,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice10_y_net
  );
  slice11 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 176,
    new_msb => 191,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice11_y_net
  );
  slice12 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 192,
    new_msb => 207,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice12_y_net
  );
  slice13 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 208,
    new_msb => 223,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice13_y_net
  );
  slice14 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 224,
    new_msb => 239,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice14_y_net
  );
  slice15 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 240,
    new_msb => 255,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice15_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/reordering extending buffer real_2/Vector Reinterpret
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_reinterpret_x8 is
  port (
    in_1 : in std_logic_vector( 16-1 downto 0 );
    in_2 : in std_logic_vector( 16-1 downto 0 );
    in_3 : in std_logic_vector( 16-1 downto 0 );
    in_4 : in std_logic_vector( 16-1 downto 0 );
    in_5 : in std_logic_vector( 16-1 downto 0 );
    in_6 : in std_logic_vector( 16-1 downto 0 );
    in_7 : in std_logic_vector( 16-1 downto 0 );
    in_8 : in std_logic_vector( 16-1 downto 0 );
    in_9 : in std_logic_vector( 16-1 downto 0 );
    in_10 : in std_logic_vector( 16-1 downto 0 );
    in_11 : in std_logic_vector( 16-1 downto 0 );
    in_12 : in std_logic_vector( 16-1 downto 0 );
    in_13 : in std_logic_vector( 16-1 downto 0 );
    in_14 : in std_logic_vector( 16-1 downto 0 );
    in_15 : in std_logic_vector( 16-1 downto 0 );
    in_16 : in std_logic_vector( 16-1 downto 0 );
    out_1 : out std_logic_vector( 16-1 downto 0 );
    out_2 : out std_logic_vector( 16-1 downto 0 );
    out_3 : out std_logic_vector( 16-1 downto 0 );
    out_4 : out std_logic_vector( 16-1 downto 0 );
    out_5 : out std_logic_vector( 16-1 downto 0 );
    out_6 : out std_logic_vector( 16-1 downto 0 );
    out_7 : out std_logic_vector( 16-1 downto 0 );
    out_8 : out std_logic_vector( 16-1 downto 0 );
    out_9 : out std_logic_vector( 16-1 downto 0 );
    out_10 : out std_logic_vector( 16-1 downto 0 );
    out_11 : out std_logic_vector( 16-1 downto 0 );
    out_12 : out std_logic_vector( 16-1 downto 0 );
    out_13 : out std_logic_vector( 16-1 downto 0 );
    out_14 : out std_logic_vector( 16-1 downto 0 );
    out_15 : out std_logic_vector( 16-1 downto 0 );
    out_16 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_vector_reinterpret_x8;
architecture structural of psb3_0_vector_reinterpret_x8 is 
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 16-1 downto 0 );
begin
  out_1 <= reinterpret0_output_port_net;
  out_2 <= reinterpret1_output_port_net;
  out_3 <= reinterpret2_output_port_net;
  out_4 <= reinterpret3_output_port_net;
  out_5 <= reinterpret4_output_port_net;
  out_6 <= reinterpret5_output_port_net;
  out_7 <= reinterpret6_output_port_net;
  out_8 <= reinterpret7_output_port_net;
  out_9 <= reinterpret8_output_port_net;
  out_10 <= reinterpret9_output_port_net;
  out_11 <= reinterpret10_output_port_net;
  out_12 <= reinterpret11_output_port_net;
  out_13 <= reinterpret12_output_port_net;
  out_14 <= reinterpret13_output_port_net;
  out_15 <= reinterpret14_output_port_net;
  out_16 <= reinterpret15_output_port_net;
  slice0_y_net <= in_1;
  slice1_y_net <= in_2;
  slice2_y_net <= in_3;
  slice3_y_net <= in_4;
  slice4_y_net <= in_5;
  slice5_y_net <= in_6;
  slice6_y_net <= in_7;
  slice7_y_net <= in_8;
  slice8_y_net <= in_9;
  slice9_y_net <= in_10;
  slice10_y_net <= in_11;
  slice11_y_net <= in_12;
  slice12_y_net <= in_13;
  slice13_y_net <= in_14;
  slice14_y_net <= in_15;
  slice15_y_net <= in_16;
  reinterpret0 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice0_y_net,
    output_port => reinterpret0_output_port_net
  );
  reinterpret1 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice1_y_net,
    output_port => reinterpret1_output_port_net
  );
  reinterpret2 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice2_y_net,
    output_port => reinterpret2_output_port_net
  );
  reinterpret3 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice3_y_net,
    output_port => reinterpret3_output_port_net
  );
  reinterpret4 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice4_y_net,
    output_port => reinterpret4_output_port_net
  );
  reinterpret5 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice5_y_net,
    output_port => reinterpret5_output_port_net
  );
  reinterpret6 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice6_y_net,
    output_port => reinterpret6_output_port_net
  );
  reinterpret7 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice7_y_net,
    output_port => reinterpret7_output_port_net
  );
  reinterpret8 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice8_y_net,
    output_port => reinterpret8_output_port_net
  );
  reinterpret9 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice9_y_net,
    output_port => reinterpret9_output_port_net
  );
  reinterpret10 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice10_y_net,
    output_port => reinterpret10_output_port_net
  );
  reinterpret11 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice11_y_net,
    output_port => reinterpret11_output_port_net
  );
  reinterpret12 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice12_y_net,
    output_port => reinterpret12_output_port_net
  );
  reinterpret13 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice13_y_net,
    output_port => reinterpret13_output_port_net
  );
  reinterpret14 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice14_y_net,
    output_port => reinterpret14_output_port_net
  );
  reinterpret15 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice15_y_net,
    output_port => reinterpret15_output_port_net
  );
end structural;
-- Generated from Simulink block PSB3_0/reordering extending buffer real_2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_reordering_extending_buffer_real_2 is
  port (
    in_reset : in std_logic_vector( 1-1 downto 0 );
    input1 : in std_logic_vector( 16-1 downto 0 );
    input2 : in std_logic_vector( 16-1 downto 0 );
    in_tvalid : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    vec_output_1 : out std_logic_vector( 16-1 downto 0 );
    vec_output_2 : out std_logic_vector( 16-1 downto 0 );
    vec_output_3 : out std_logic_vector( 16-1 downto 0 );
    vec_output_4 : out std_logic_vector( 16-1 downto 0 );
    vec_output_5 : out std_logic_vector( 16-1 downto 0 );
    vec_output_6 : out std_logic_vector( 16-1 downto 0 );
    vec_output_7 : out std_logic_vector( 16-1 downto 0 );
    vec_output_8 : out std_logic_vector( 16-1 downto 0 );
    vec_output_9 : out std_logic_vector( 16-1 downto 0 );
    vec_output_10 : out std_logic_vector( 16-1 downto 0 );
    vec_output_11 : out std_logic_vector( 16-1 downto 0 );
    vec_output_12 : out std_logic_vector( 16-1 downto 0 );
    vec_output_13 : out std_logic_vector( 16-1 downto 0 );
    vec_output_14 : out std_logic_vector( 16-1 downto 0 );
    vec_output_15 : out std_logic_vector( 16-1 downto 0 );
    vec_output_16 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_reordering_extending_buffer_real_2;
architecture structural of psb3_0_reordering_extending_buffer_real_2 is 
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal delay19_q_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal slice3_y_net : std_logic_vector( 16-1 downto 0 );
  signal ce_net : std_logic;
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mux1_y_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal gin_tl_reset_net : std_logic_vector( 1-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 16-1 downto 0 );
  signal mux5_y_net_x0 : std_logic_vector( 256-1 downto 0 );
  signal mux5_y_net : std_logic_vector( 16-1 downto 0 );
  signal bitbasher1_out_x0_net : std_logic_vector( 256-1 downto 0 );
  signal dual_port_ram_1_douta_net : std_logic_vector( 16-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 1-1 downto 0 );
  signal delay10_q_net : std_logic_vector( 1-1 downto 0 );
  signal single_port_ram_data_out_net : std_logic_vector( 1-1 downto 0 );
  signal dual_port_ram_1_doutb_net : std_logic_vector( 16-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 16-1 downto 0 );
  signal delay11_q_net : std_logic_vector( 1-1 downto 0 );
  signal we_0 : std_logic_vector( 1-1 downto 0 );
  signal dual_port_ram_0_doutb_net : std_logic_vector( 16-1 downto 0 );
  signal dual_port_ram_0_douta_net : std_logic_vector( 16-1 downto 0 );
  signal constant2_op_net : std_logic_vector( 1-1 downto 0 );
  signal bitbasher_out_x0_net : std_logic_vector( 256-1 downto 0 );
  signal constant_op_net : std_logic_vector( 1-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 9-1 downto 0 );
  signal delay7_q_net : std_logic_vector( 8-1 downto 0 );
  signal delay9_q_net : std_logic_vector( 1-1 downto 0 );
  signal inverter_op_net : std_logic_vector( 1-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 1-1 downto 0 );
  signal even_addr_w_op_net : std_logic_vector( 9-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 16-1 downto 0 );
  signal addr_r_op_net : std_logic_vector( 8-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 9-1 downto 0 );
  signal odd_addr_w_op_net : std_logic_vector( 9-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux4_y_net : std_logic_vector( 9-1 downto 0 );
  signal out_in_1024_out_x0_net : std_logic_vector( 9-1 downto 0 );
  signal mux3_y_net : std_logic_vector( 9-1 downto 0 );
  signal mux2_y_net : std_logic_vector( 9-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 9-1 downto 0 );
  signal addr_control_op_net : std_logic_vector( 9-1 downto 0 );
begin
  vec_output_1 <= reinterpret0_output_port_net;
  vec_output_2 <= reinterpret1_output_port_net;
  vec_output_3 <= reinterpret2_output_port_net;
  vec_output_4 <= reinterpret3_output_port_net;
  vec_output_5 <= reinterpret4_output_port_net;
  vec_output_6 <= reinterpret5_output_port_net;
  vec_output_7 <= reinterpret6_output_port_net;
  vec_output_8 <= reinterpret7_output_port_net;
  vec_output_9 <= reinterpret8_output_port_net;
  vec_output_10 <= reinterpret9_output_port_net;
  vec_output_11 <= reinterpret10_output_port_net;
  vec_output_12 <= reinterpret11_output_port_net;
  vec_output_13 <= reinterpret12_output_port_net;
  vec_output_14 <= reinterpret13_output_port_net;
  vec_output_15 <= reinterpret14_output_port_net;
  vec_output_16 <= reinterpret15_output_port_net;
  gin_tl_reset_net <= in_reset;
  mux1_y_net_x0 <= input1;
  mux5_y_net <= input2;
  delay19_q_net <= in_tvalid;
  clk_net <= clk_1;
  ce_net <= ce_1;
  scalar_to_vector4 : entity xil_defaultlib.psb3_0_scalar_to_vector4_x5 
  port map (
    i => mux5_y_net_x0,
    o_1 => slice0_y_net,
    o_2 => slice1_y_net,
    o_3 => slice2_y_net,
    o_4 => slice3_y_net,
    o_5 => slice4_y_net,
    o_6 => slice5_y_net,
    o_7 => slice6_y_net,
    o_8 => slice7_y_net,
    o_9 => slice8_y_net,
    o_10 => slice9_y_net,
    o_11 => slice10_y_net,
    o_12 => slice11_y_net,
    o_13 => slice12_y_net,
    o_14 => slice13_y_net,
    o_15 => slice14_y_net,
    o_16 => slice15_y_net
  );
  vector_reinterpret : entity xil_defaultlib.psb3_0_vector_reinterpret_x8 
  port map (
    in_1 => slice0_y_net,
    in_2 => slice1_y_net,
    in_3 => slice2_y_net,
    in_4 => slice3_y_net,
    in_5 => slice4_y_net,
    in_6 => slice5_y_net,
    in_7 => slice6_y_net,
    in_8 => slice7_y_net,
    in_9 => slice8_y_net,
    in_10 => slice9_y_net,
    in_11 => slice10_y_net,
    in_12 => slice11_y_net,
    in_13 => slice12_y_net,
    in_14 => slice13_y_net,
    in_15 => slice14_y_net,
    in_16 => slice15_y_net,
    out_1 => reinterpret0_output_port_net,
    out_2 => reinterpret1_output_port_net,
    out_3 => reinterpret2_output_port_net,
    out_4 => reinterpret3_output_port_net,
    out_5 => reinterpret4_output_port_net,
    out_6 => reinterpret5_output_port_net,
    out_7 => reinterpret6_output_port_net,
    out_8 => reinterpret7_output_port_net,
    out_9 => reinterpret8_output_port_net,
    out_10 => reinterpret9_output_port_net,
    out_11 => reinterpret10_output_port_net,
    out_12 => reinterpret11_output_port_net,
    out_13 => reinterpret12_output_port_net,
    out_14 => reinterpret13_output_port_net,
    out_15 => reinterpret14_output_port_net,
    out_16 => reinterpret15_output_port_net
  );
  bitbasher : entity xil_defaultlib.sysgen_bitbasher_4648460ba6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    a => dual_port_ram_0_douta_net,
    b => dual_port_ram_0_doutb_net,
    out_x0 => bitbasher_out_x0_net
  );
  bitbasher1 : entity xil_defaultlib.sysgen_bitbasher_4648460ba6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    a => dual_port_ram_1_douta_net,
    b => dual_port_ram_1_doutb_net,
    out_x0 => bitbasher1_out_x0_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_de9059c03f 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_71e89d757c 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  constant2 : entity xil_defaultlib.sysgen_constant_71e89d757c 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant2_op_net
  );
  delay : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => single_port_ram_data_out_net,
    clk => clk_net,
    ce => ce_net,
    q => we_0
  );
  delay1 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 16
  )
  port map (
    en => '1',
    rst => '0',
    d => mux1_y_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay10 : entity xil_defaultlib.sysgen_delay_906db00812 
  port map (
    clr => '0',
    d => constant1_op_net,
    rst => gin_tl_reset_net,
    clk => clk_net,
    ce => ce_net,
    q => delay10_q_net
  );
  delay11 : entity xil_defaultlib.sysgen_delay_906db00812 
  port map (
    clr => '0',
    d => constant2_op_net,
    rst => gin_tl_reset_net,
    clk => clk_net,
    ce => ce_net,
    q => delay11_q_net
  );
  delay2 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 16
  )
  port map (
    en => '1',
    rst => '0',
    d => mux5_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay3 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => we_0,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  delay4 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => inverter_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net
  );
  delay5 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 9
  )
  port map (
    en => '1',
    rst => '0',
    d => even_addr_w_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  delay6 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 9
  )
  port map (
    en => '1',
    rst => '0',
    d => odd_addr_w_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay6_q_net
  );
  delay7 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 8
  )
  port map (
    en => '1',
    rst => '0',
    d => addr_r_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay7_q_net
  );
  delay9 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay9_q_net
  );
  dual_port_ram_0 : entity xil_defaultlib.psb3_0_xltdpram 
  generic map (
    addr_width_b => 9,
    clocking_mode => "common_clock",
    data_width_b => 16,
    latency => 1,
    mem_init_file => "xpm_c5fd30_vivado.mem",
    mem_size => 8192,
    mem_type => "block",
    read_reset_a => "0",
    read_reset_b => "0",
    width => 16,
    width_addr => 9,
    write_mode_a => "read_first",
    write_mode_b => "read_first"
  )
  port map (
    ena => "1",
    rsta => "0",
    rstb => "0",
    addra => mux1_y_net,
    dina => delay1_q_net,
    wea => delay3_q_net,
    addrb => mux2_y_net,
    dinb => delay2_q_net,
    web => delay3_q_net,
    enb => delay11_q_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dual_port_ram_0_douta_net,
    doutb => dual_port_ram_0_doutb_net
  );
  dual_port_ram_1 : entity xil_defaultlib.psb3_0_xltdpram 
  generic map (
    addr_width_b => 9,
    clocking_mode => "common_clock",
    data_width_b => 16,
    latency => 1,
    mem_init_file => "xpm_c5fd30_vivado.mem",
    mem_size => 8192,
    mem_type => "block",
    read_reset_a => "0",
    read_reset_b => "0",
    width => 16,
    width_addr => 9,
    write_mode_a => "read_first",
    write_mode_b => "read_first"
  )
  port map (
    ena => "1",
    rsta => "0",
    rstb => "0",
    addra => mux3_y_net,
    dina => delay1_q_net,
    wea => delay4_q_net,
    addrb => mux4_y_net,
    dinb => delay2_q_net,
    web => delay4_q_net,
    enb => delay10_q_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dual_port_ram_1_douta_net,
    doutb => dual_port_ram_1_doutb_net
  );
  inverter : entity xil_defaultlib.sysgen_inverter_ac5174c184 
  port map (
    clr => '0',
    ip => single_port_ram_data_out_net,
    clk => clk_net,
    ce => ce_net,
    op => inverter_op_net
  );
  mux1 : entity xil_defaultlib.sysgen_mux_303302b1e4 
  port map (
    clr => '0',
    sel => we_0,
    d0 => delay7_q_net,
    d1 => delay5_q_net,
    clk => clk_net,
    ce => ce_net,
    y => mux1_y_net
  );
  mux2 : entity xil_defaultlib.sysgen_mux_c7d0cfa098 
  port map (
    clr => '0',
    sel => we_0,
    d0 => out_in_1024_out_x0_net,
    d1 => delay6_q_net,
    clk => clk_net,
    ce => ce_net,
    y => mux2_y_net
  );
  mux3 : entity xil_defaultlib.sysgen_mux_303302b1e4 
  port map (
    clr => '0',
    sel => inverter_op_net,
    d0 => delay7_q_net,
    d1 => delay5_q_net,
    clk => clk_net,
    ce => ce_net,
    y => mux3_y_net
  );
  mux4 : entity xil_defaultlib.sysgen_mux_c7d0cfa098 
  port map (
    clr => '0',
    sel => inverter_op_net,
    d0 => out_in_1024_out_x0_net,
    d1 => delay6_q_net,
    clk => clk_net,
    ce => ce_net,
    y => mux4_y_net
  );
  mux5 : entity xil_defaultlib.sysgen_mux_1f606cf16b 
  port map (
    clr => '0',
    sel => delay9_q_net,
    d0 => bitbasher_out_x0_net,
    d1 => bitbasher1_out_x0_net,
    clk => clk_net,
    ce => ce_net,
    y => mux5_y_net_x0
  );
  single_port_ram : entity xil_defaultlib.psb3_0_xlspram 
  generic map (
    init_value => b"0",
    latency => 1,
    mem_init_file => "xpm_95b604_vivado.mem",
    mem_size => 512,
    mem_type => "block",
    read_reset_val => "0",
    width => 1,
    width_addr => 9,
    write_mode_a => "read_first",
    xpm_lat => 1
  )
  port map (
    en => "1",
    rst => "0",
    addr => addr_control_op_net,
    data_in => constant_op_net,
    we => constant_op_net,
    clk => clk_net,
    ce => ce_net,
    data_out => single_port_ram_data_out_net
  );
  addr_control : entity xil_defaultlib.psb3_0_xlcounter_free 
  generic map (
    core_name0 => "psb3_0_c_counter_binary_v12_0_i4",
    op_arith => xlUnsigned,
    op_width => 9
  )
  port map (
    clr => '0',
    rst => gin_tl_reset_net,
    en => delay19_q_net,
    clk => clk_net,
    ce => ce_net,
    op => addr_control_op_net
  );
  addr_r : entity xil_defaultlib.psb3_0_xlcounter_free 
  generic map (
    core_name0 => "psb3_0_c_counter_binary_v12_0_i3",
    op_arith => xlUnsigned,
    op_width => 8
  )
  port map (
    clr => '0',
    rst => gin_tl_reset_net,
    en => delay19_q_net,
    clk => clk_net,
    ce => ce_net,
    op => addr_r_op_net
  );
  even_addr_w : entity xil_defaultlib.psb3_0_xlcounter_free 
  generic map (
    core_name0 => "psb3_0_c_counter_binary_v12_0_i5",
    op_arith => xlUnsigned,
    op_width => 9
  )
  port map (
    clr => '0',
    rst => gin_tl_reset_net,
    en => delay19_q_net,
    clk => clk_net,
    ce => ce_net,
    op => even_addr_w_op_net
  );
  odd_addr_w : entity xil_defaultlib.psb3_0_xlcounter_free 
  generic map (
    core_name0 => "psb3_0_c_counter_binary_v12_0_i6",
    op_arith => xlUnsigned,
    op_width => 9
  )
  port map (
    clr => '0',
    rst => gin_tl_reset_net,
    en => delay19_q_net,
    clk => clk_net,
    ce => ce_net,
    op => odd_addr_w_op_net
  );
  out_in_1024 : entity xil_defaultlib.sysgen_bitbasher_a62d2ce679 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in_x0 => delay7_q_net,
    out_x0 => out_in_1024_out_x0_net
  );
end structural;
-- Generated from Simulink block PSB3_0/reordering extending buffer real_3/Scalar to Vector4
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_scalar_to_vector4_x6 is
  port (
    i : in std_logic_vector( 256-1 downto 0 );
    o_1 : out std_logic_vector( 16-1 downto 0 );
    o_2 : out std_logic_vector( 16-1 downto 0 );
    o_3 : out std_logic_vector( 16-1 downto 0 );
    o_4 : out std_logic_vector( 16-1 downto 0 );
    o_5 : out std_logic_vector( 16-1 downto 0 );
    o_6 : out std_logic_vector( 16-1 downto 0 );
    o_7 : out std_logic_vector( 16-1 downto 0 );
    o_8 : out std_logic_vector( 16-1 downto 0 );
    o_9 : out std_logic_vector( 16-1 downto 0 );
    o_10 : out std_logic_vector( 16-1 downto 0 );
    o_11 : out std_logic_vector( 16-1 downto 0 );
    o_12 : out std_logic_vector( 16-1 downto 0 );
    o_13 : out std_logic_vector( 16-1 downto 0 );
    o_14 : out std_logic_vector( 16-1 downto 0 );
    o_15 : out std_logic_vector( 16-1 downto 0 );
    o_16 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_scalar_to_vector4_x6;
architecture structural of psb3_0_scalar_to_vector4_x6 is 
  signal slice9_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 16-1 downto 0 );
  signal mux5_y_net : std_logic_vector( 256-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 16-1 downto 0 );
begin
  o_1 <= slice0_y_net;
  o_2 <= slice1_y_net;
  o_3 <= slice2_y_net;
  o_4 <= slice3_y_net;
  o_5 <= slice4_y_net;
  o_6 <= slice5_y_net;
  o_7 <= slice6_y_net;
  o_8 <= slice7_y_net;
  o_9 <= slice8_y_net;
  o_10 <= slice9_y_net;
  o_11 <= slice10_y_net;
  o_12 <= slice11_y_net;
  o_13 <= slice12_y_net;
  o_14 <= slice13_y_net;
  o_15 <= slice14_y_net;
  o_16 <= slice15_y_net;
  mux5_y_net <= i;
  slice0 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 15,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice0_y_net
  );
  slice1 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 16,
    new_msb => 31,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice1_y_net
  );
  slice2 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 32,
    new_msb => 47,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice2_y_net
  );
  slice3 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 48,
    new_msb => 63,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice3_y_net
  );
  slice4 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 64,
    new_msb => 79,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice4_y_net
  );
  slice5 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 80,
    new_msb => 95,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice5_y_net
  );
  slice6 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 96,
    new_msb => 111,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice6_y_net
  );
  slice7 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 112,
    new_msb => 127,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice7_y_net
  );
  slice8 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 128,
    new_msb => 143,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice8_y_net
  );
  slice9 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 144,
    new_msb => 159,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice9_y_net
  );
  slice10 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 160,
    new_msb => 175,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice10_y_net
  );
  slice11 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 176,
    new_msb => 191,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice11_y_net
  );
  slice12 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 192,
    new_msb => 207,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice12_y_net
  );
  slice13 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 208,
    new_msb => 223,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice13_y_net
  );
  slice14 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 224,
    new_msb => 239,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice14_y_net
  );
  slice15 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 240,
    new_msb => 255,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice15_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/reordering extending buffer real_3/Vector Reinterpret
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_reinterpret_x9 is
  port (
    in_1 : in std_logic_vector( 16-1 downto 0 );
    in_2 : in std_logic_vector( 16-1 downto 0 );
    in_3 : in std_logic_vector( 16-1 downto 0 );
    in_4 : in std_logic_vector( 16-1 downto 0 );
    in_5 : in std_logic_vector( 16-1 downto 0 );
    in_6 : in std_logic_vector( 16-1 downto 0 );
    in_7 : in std_logic_vector( 16-1 downto 0 );
    in_8 : in std_logic_vector( 16-1 downto 0 );
    in_9 : in std_logic_vector( 16-1 downto 0 );
    in_10 : in std_logic_vector( 16-1 downto 0 );
    in_11 : in std_logic_vector( 16-1 downto 0 );
    in_12 : in std_logic_vector( 16-1 downto 0 );
    in_13 : in std_logic_vector( 16-1 downto 0 );
    in_14 : in std_logic_vector( 16-1 downto 0 );
    in_15 : in std_logic_vector( 16-1 downto 0 );
    in_16 : in std_logic_vector( 16-1 downto 0 );
    out_1 : out std_logic_vector( 16-1 downto 0 );
    out_2 : out std_logic_vector( 16-1 downto 0 );
    out_3 : out std_logic_vector( 16-1 downto 0 );
    out_4 : out std_logic_vector( 16-1 downto 0 );
    out_5 : out std_logic_vector( 16-1 downto 0 );
    out_6 : out std_logic_vector( 16-1 downto 0 );
    out_7 : out std_logic_vector( 16-1 downto 0 );
    out_8 : out std_logic_vector( 16-1 downto 0 );
    out_9 : out std_logic_vector( 16-1 downto 0 );
    out_10 : out std_logic_vector( 16-1 downto 0 );
    out_11 : out std_logic_vector( 16-1 downto 0 );
    out_12 : out std_logic_vector( 16-1 downto 0 );
    out_13 : out std_logic_vector( 16-1 downto 0 );
    out_14 : out std_logic_vector( 16-1 downto 0 );
    out_15 : out std_logic_vector( 16-1 downto 0 );
    out_16 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_vector_reinterpret_x9;
architecture structural of psb3_0_vector_reinterpret_x9 is 
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 16-1 downto 0 );
begin
  out_1 <= reinterpret0_output_port_net;
  out_2 <= reinterpret1_output_port_net;
  out_3 <= reinterpret2_output_port_net;
  out_4 <= reinterpret3_output_port_net;
  out_5 <= reinterpret4_output_port_net;
  out_6 <= reinterpret5_output_port_net;
  out_7 <= reinterpret6_output_port_net;
  out_8 <= reinterpret7_output_port_net;
  out_9 <= reinterpret8_output_port_net;
  out_10 <= reinterpret9_output_port_net;
  out_11 <= reinterpret10_output_port_net;
  out_12 <= reinterpret11_output_port_net;
  out_13 <= reinterpret12_output_port_net;
  out_14 <= reinterpret13_output_port_net;
  out_15 <= reinterpret14_output_port_net;
  out_16 <= reinterpret15_output_port_net;
  slice0_y_net <= in_1;
  slice1_y_net <= in_2;
  slice2_y_net <= in_3;
  slice3_y_net <= in_4;
  slice4_y_net <= in_5;
  slice5_y_net <= in_6;
  slice6_y_net <= in_7;
  slice7_y_net <= in_8;
  slice8_y_net <= in_9;
  slice9_y_net <= in_10;
  slice10_y_net <= in_11;
  slice11_y_net <= in_12;
  slice12_y_net <= in_13;
  slice13_y_net <= in_14;
  slice14_y_net <= in_15;
  slice15_y_net <= in_16;
  reinterpret0 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice0_y_net,
    output_port => reinterpret0_output_port_net
  );
  reinterpret1 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice1_y_net,
    output_port => reinterpret1_output_port_net
  );
  reinterpret2 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice2_y_net,
    output_port => reinterpret2_output_port_net
  );
  reinterpret3 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice3_y_net,
    output_port => reinterpret3_output_port_net
  );
  reinterpret4 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice4_y_net,
    output_port => reinterpret4_output_port_net
  );
  reinterpret5 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice5_y_net,
    output_port => reinterpret5_output_port_net
  );
  reinterpret6 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice6_y_net,
    output_port => reinterpret6_output_port_net
  );
  reinterpret7 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice7_y_net,
    output_port => reinterpret7_output_port_net
  );
  reinterpret8 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice8_y_net,
    output_port => reinterpret8_output_port_net
  );
  reinterpret9 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice9_y_net,
    output_port => reinterpret9_output_port_net
  );
  reinterpret10 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice10_y_net,
    output_port => reinterpret10_output_port_net
  );
  reinterpret11 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice11_y_net,
    output_port => reinterpret11_output_port_net
  );
  reinterpret12 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice12_y_net,
    output_port => reinterpret12_output_port_net
  );
  reinterpret13 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice13_y_net,
    output_port => reinterpret13_output_port_net
  );
  reinterpret14 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice14_y_net,
    output_port => reinterpret14_output_port_net
  );
  reinterpret15 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice15_y_net,
    output_port => reinterpret15_output_port_net
  );
end structural;
-- Generated from Simulink block PSB3_0/reordering extending buffer real_3
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_reordering_extending_buffer_real_3 is
  port (
    in_reset : in std_logic_vector( 1-1 downto 0 );
    input1 : in std_logic_vector( 16-1 downto 0 );
    input2 : in std_logic_vector( 16-1 downto 0 );
    in_tvalid : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    vec_output_1 : out std_logic_vector( 16-1 downto 0 );
    vec_output_2 : out std_logic_vector( 16-1 downto 0 );
    vec_output_3 : out std_logic_vector( 16-1 downto 0 );
    vec_output_4 : out std_logic_vector( 16-1 downto 0 );
    vec_output_5 : out std_logic_vector( 16-1 downto 0 );
    vec_output_6 : out std_logic_vector( 16-1 downto 0 );
    vec_output_7 : out std_logic_vector( 16-1 downto 0 );
    vec_output_8 : out std_logic_vector( 16-1 downto 0 );
    vec_output_9 : out std_logic_vector( 16-1 downto 0 );
    vec_output_10 : out std_logic_vector( 16-1 downto 0 );
    vec_output_11 : out std_logic_vector( 16-1 downto 0 );
    vec_output_12 : out std_logic_vector( 16-1 downto 0 );
    vec_output_13 : out std_logic_vector( 16-1 downto 0 );
    vec_output_14 : out std_logic_vector( 16-1 downto 0 );
    vec_output_15 : out std_logic_vector( 16-1 downto 0 );
    vec_output_16 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_reordering_extending_buffer_real_3;
architecture structural of psb3_0_reordering_extending_buffer_real_3 is 
  signal delay3_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 9-1 downto 0 );
  signal mux2_y_net : std_logic_vector( 9-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 9-1 downto 0 );
  signal delay7_q_net : std_logic_vector( 8-1 downto 0 );
  signal inverter_op_net : std_logic_vector( 1-1 downto 0 );
  signal delay9_q_net : std_logic_vector( 1-1 downto 0 );
  signal even_addr_w_op_net : std_logic_vector( 9-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 9-1 downto 0 );
  signal odd_addr_w_op_net : std_logic_vector( 9-1 downto 0 );
  signal addr_r_op_net : std_logic_vector( 8-1 downto 0 );
  signal mux4_y_net : std_logic_vector( 9-1 downto 0 );
  signal addr_control_op_net : std_logic_vector( 9-1 downto 0 );
  signal mux3_y_net : std_logic_vector( 9-1 downto 0 );
  signal out_in_1024_out_x0_net : std_logic_vector( 9-1 downto 0 );
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 16-1 downto 0 );
  signal dual_port_ram_0_doutb_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal ce_net : std_logic;
  signal mux2_y_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal bitbasher_out_x0_net : std_logic_vector( 256-1 downto 0 );
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 16-1 downto 0 );
  signal gin_tl_reset_net : std_logic_vector( 1-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 16-1 downto 0 );
  signal mux5_y_net : std_logic_vector( 256-1 downto 0 );
  signal dual_port_ram_0_douta_net : std_logic_vector( 16-1 downto 0 );
  signal delay19_q_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal clk_net : std_logic;
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mux6_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 16-1 downto 0 );
  signal delay11_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 16-1 downto 0 );
  signal constant_op_net : std_logic_vector( 1-1 downto 0 );
  signal single_port_ram_data_out_net : std_logic_vector( 1-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 16-1 downto 0 );
  signal dual_port_ram_1_douta_net : std_logic_vector( 16-1 downto 0 );
  signal we_0 : std_logic_vector( 1-1 downto 0 );
  signal dual_port_ram_1_doutb_net : std_logic_vector( 16-1 downto 0 );
  signal bitbasher1_out_x0_net : std_logic_vector( 256-1 downto 0 );
  signal constant2_op_net : std_logic_vector( 1-1 downto 0 );
  signal delay10_q_net : std_logic_vector( 1-1 downto 0 );
begin
  vec_output_1 <= reinterpret0_output_port_net;
  vec_output_2 <= reinterpret1_output_port_net;
  vec_output_3 <= reinterpret2_output_port_net;
  vec_output_4 <= reinterpret3_output_port_net;
  vec_output_5 <= reinterpret4_output_port_net;
  vec_output_6 <= reinterpret5_output_port_net;
  vec_output_7 <= reinterpret6_output_port_net;
  vec_output_8 <= reinterpret7_output_port_net;
  vec_output_9 <= reinterpret8_output_port_net;
  vec_output_10 <= reinterpret9_output_port_net;
  vec_output_11 <= reinterpret10_output_port_net;
  vec_output_12 <= reinterpret11_output_port_net;
  vec_output_13 <= reinterpret12_output_port_net;
  vec_output_14 <= reinterpret13_output_port_net;
  vec_output_15 <= reinterpret14_output_port_net;
  vec_output_16 <= reinterpret15_output_port_net;
  gin_tl_reset_net <= in_reset;
  mux2_y_net_x0 <= input1;
  mux6_y_net <= input2;
  delay19_q_net <= in_tvalid;
  clk_net <= clk_1;
  ce_net <= ce_1;
  scalar_to_vector4 : entity xil_defaultlib.psb3_0_scalar_to_vector4_x6 
  port map (
    i => mux5_y_net,
    o_1 => slice0_y_net,
    o_2 => slice1_y_net,
    o_3 => slice2_y_net,
    o_4 => slice3_y_net,
    o_5 => slice4_y_net,
    o_6 => slice5_y_net,
    o_7 => slice6_y_net,
    o_8 => slice7_y_net,
    o_9 => slice8_y_net,
    o_10 => slice9_y_net,
    o_11 => slice10_y_net,
    o_12 => slice11_y_net,
    o_13 => slice12_y_net,
    o_14 => slice13_y_net,
    o_15 => slice14_y_net,
    o_16 => slice15_y_net
  );
  vector_reinterpret : entity xil_defaultlib.psb3_0_vector_reinterpret_x9 
  port map (
    in_1 => slice0_y_net,
    in_2 => slice1_y_net,
    in_3 => slice2_y_net,
    in_4 => slice3_y_net,
    in_5 => slice4_y_net,
    in_6 => slice5_y_net,
    in_7 => slice6_y_net,
    in_8 => slice7_y_net,
    in_9 => slice8_y_net,
    in_10 => slice9_y_net,
    in_11 => slice10_y_net,
    in_12 => slice11_y_net,
    in_13 => slice12_y_net,
    in_14 => slice13_y_net,
    in_15 => slice14_y_net,
    in_16 => slice15_y_net,
    out_1 => reinterpret0_output_port_net,
    out_2 => reinterpret1_output_port_net,
    out_3 => reinterpret2_output_port_net,
    out_4 => reinterpret3_output_port_net,
    out_5 => reinterpret4_output_port_net,
    out_6 => reinterpret5_output_port_net,
    out_7 => reinterpret6_output_port_net,
    out_8 => reinterpret7_output_port_net,
    out_9 => reinterpret8_output_port_net,
    out_10 => reinterpret9_output_port_net,
    out_11 => reinterpret10_output_port_net,
    out_12 => reinterpret11_output_port_net,
    out_13 => reinterpret12_output_port_net,
    out_14 => reinterpret13_output_port_net,
    out_15 => reinterpret14_output_port_net,
    out_16 => reinterpret15_output_port_net
  );
  bitbasher : entity xil_defaultlib.sysgen_bitbasher_4648460ba6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    a => dual_port_ram_0_douta_net,
    b => dual_port_ram_0_doutb_net,
    out_x0 => bitbasher_out_x0_net
  );
  bitbasher1 : entity xil_defaultlib.sysgen_bitbasher_4648460ba6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    a => dual_port_ram_1_douta_net,
    b => dual_port_ram_1_doutb_net,
    out_x0 => bitbasher1_out_x0_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_de9059c03f 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_71e89d757c 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  constant2 : entity xil_defaultlib.sysgen_constant_71e89d757c 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant2_op_net
  );
  delay : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => single_port_ram_data_out_net,
    clk => clk_net,
    ce => ce_net,
    q => we_0
  );
  delay1 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 16
  )
  port map (
    en => '1',
    rst => '0',
    d => mux2_y_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay10 : entity xil_defaultlib.sysgen_delay_906db00812 
  port map (
    clr => '0',
    d => constant1_op_net,
    rst => gin_tl_reset_net,
    clk => clk_net,
    ce => ce_net,
    q => delay10_q_net
  );
  delay11 : entity xil_defaultlib.sysgen_delay_906db00812 
  port map (
    clr => '0',
    d => constant2_op_net,
    rst => gin_tl_reset_net,
    clk => clk_net,
    ce => ce_net,
    q => delay11_q_net
  );
  delay2 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 16
  )
  port map (
    en => '1',
    rst => '0',
    d => mux6_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay3 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => we_0,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  delay4 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => inverter_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net
  );
  delay5 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 9
  )
  port map (
    en => '1',
    rst => '0',
    d => even_addr_w_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  delay6 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 9
  )
  port map (
    en => '1',
    rst => '0',
    d => odd_addr_w_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay6_q_net
  );
  delay7 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 8
  )
  port map (
    en => '1',
    rst => '0',
    d => addr_r_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay7_q_net
  );
  delay9 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay9_q_net
  );
  dual_port_ram_0 : entity xil_defaultlib.psb3_0_xltdpram 
  generic map (
    addr_width_b => 9,
    clocking_mode => "common_clock",
    data_width_b => 16,
    latency => 1,
    mem_init_file => "xpm_c5fd30_vivado.mem",
    mem_size => 8192,
    mem_type => "block",
    read_reset_a => "0",
    read_reset_b => "0",
    width => 16,
    width_addr => 9,
    write_mode_a => "read_first",
    write_mode_b => "read_first"
  )
  port map (
    ena => "1",
    rsta => "0",
    rstb => "0",
    addra => mux1_y_net,
    dina => delay1_q_net,
    wea => delay3_q_net,
    addrb => mux2_y_net,
    dinb => delay2_q_net,
    web => delay3_q_net,
    enb => delay11_q_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dual_port_ram_0_douta_net,
    doutb => dual_port_ram_0_doutb_net
  );
  dual_port_ram_1 : entity xil_defaultlib.psb3_0_xltdpram 
  generic map (
    addr_width_b => 9,
    clocking_mode => "common_clock",
    data_width_b => 16,
    latency => 1,
    mem_init_file => "xpm_c5fd30_vivado.mem",
    mem_size => 8192,
    mem_type => "block",
    read_reset_a => "0",
    read_reset_b => "0",
    width => 16,
    width_addr => 9,
    write_mode_a => "read_first",
    write_mode_b => "read_first"
  )
  port map (
    ena => "1",
    rsta => "0",
    rstb => "0",
    addra => mux3_y_net,
    dina => delay1_q_net,
    wea => delay4_q_net,
    addrb => mux4_y_net,
    dinb => delay2_q_net,
    web => delay4_q_net,
    enb => delay10_q_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dual_port_ram_1_douta_net,
    doutb => dual_port_ram_1_doutb_net
  );
  inverter : entity xil_defaultlib.sysgen_inverter_ac5174c184 
  port map (
    clr => '0',
    ip => single_port_ram_data_out_net,
    clk => clk_net,
    ce => ce_net,
    op => inverter_op_net
  );
  mux1 : entity xil_defaultlib.sysgen_mux_303302b1e4 
  port map (
    clr => '0',
    sel => we_0,
    d0 => delay7_q_net,
    d1 => delay5_q_net,
    clk => clk_net,
    ce => ce_net,
    y => mux1_y_net
  );
  mux2 : entity xil_defaultlib.sysgen_mux_c7d0cfa098 
  port map (
    clr => '0',
    sel => we_0,
    d0 => out_in_1024_out_x0_net,
    d1 => delay6_q_net,
    clk => clk_net,
    ce => ce_net,
    y => mux2_y_net
  );
  mux3 : entity xil_defaultlib.sysgen_mux_303302b1e4 
  port map (
    clr => '0',
    sel => inverter_op_net,
    d0 => delay7_q_net,
    d1 => delay5_q_net,
    clk => clk_net,
    ce => ce_net,
    y => mux3_y_net
  );
  mux4 : entity xil_defaultlib.sysgen_mux_c7d0cfa098 
  port map (
    clr => '0',
    sel => inverter_op_net,
    d0 => out_in_1024_out_x0_net,
    d1 => delay6_q_net,
    clk => clk_net,
    ce => ce_net,
    y => mux4_y_net
  );
  mux5 : entity xil_defaultlib.sysgen_mux_1f606cf16b 
  port map (
    clr => '0',
    sel => delay9_q_net,
    d0 => bitbasher_out_x0_net,
    d1 => bitbasher1_out_x0_net,
    clk => clk_net,
    ce => ce_net,
    y => mux5_y_net
  );
  single_port_ram : entity xil_defaultlib.psb3_0_xlspram 
  generic map (
    init_value => b"0",
    latency => 1,
    mem_init_file => "xpm_95b604_vivado.mem",
    mem_size => 512,
    mem_type => "block",
    read_reset_val => "0",
    width => 1,
    width_addr => 9,
    write_mode_a => "read_first",
    xpm_lat => 1
  )
  port map (
    en => "1",
    rst => "0",
    addr => addr_control_op_net,
    data_in => constant_op_net,
    we => constant_op_net,
    clk => clk_net,
    ce => ce_net,
    data_out => single_port_ram_data_out_net
  );
  addr_control : entity xil_defaultlib.psb3_0_xlcounter_free 
  generic map (
    core_name0 => "psb3_0_c_counter_binary_v12_0_i4",
    op_arith => xlUnsigned,
    op_width => 9
  )
  port map (
    clr => '0',
    rst => gin_tl_reset_net,
    en => delay19_q_net,
    clk => clk_net,
    ce => ce_net,
    op => addr_control_op_net
  );
  addr_r : entity xil_defaultlib.psb3_0_xlcounter_free 
  generic map (
    core_name0 => "psb3_0_c_counter_binary_v12_0_i3",
    op_arith => xlUnsigned,
    op_width => 8
  )
  port map (
    clr => '0',
    rst => gin_tl_reset_net,
    en => delay19_q_net,
    clk => clk_net,
    ce => ce_net,
    op => addr_r_op_net
  );
  even_addr_w : entity xil_defaultlib.psb3_0_xlcounter_free 
  generic map (
    core_name0 => "psb3_0_c_counter_binary_v12_0_i5",
    op_arith => xlUnsigned,
    op_width => 9
  )
  port map (
    clr => '0',
    rst => gin_tl_reset_net,
    en => delay19_q_net,
    clk => clk_net,
    ce => ce_net,
    op => even_addr_w_op_net
  );
  odd_addr_w : entity xil_defaultlib.psb3_0_xlcounter_free 
  generic map (
    core_name0 => "psb3_0_c_counter_binary_v12_0_i6",
    op_arith => xlUnsigned,
    op_width => 9
  )
  port map (
    clr => '0',
    rst => gin_tl_reset_net,
    en => delay19_q_net,
    clk => clk_net,
    ce => ce_net,
    op => odd_addr_w_op_net
  );
  out_in_1024 : entity xil_defaultlib.sysgen_bitbasher_a62d2ce679 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in_x0 => delay7_q_net,
    out_x0 => out_in_1024_out_x0_net
  );
end structural;
-- Generated from Simulink block PSB3_0/reordering extending buffer real_4/Scalar to Vector4
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_scalar_to_vector4_x7 is
  port (
    i : in std_logic_vector( 256-1 downto 0 );
    o_1 : out std_logic_vector( 16-1 downto 0 );
    o_2 : out std_logic_vector( 16-1 downto 0 );
    o_3 : out std_logic_vector( 16-1 downto 0 );
    o_4 : out std_logic_vector( 16-1 downto 0 );
    o_5 : out std_logic_vector( 16-1 downto 0 );
    o_6 : out std_logic_vector( 16-1 downto 0 );
    o_7 : out std_logic_vector( 16-1 downto 0 );
    o_8 : out std_logic_vector( 16-1 downto 0 );
    o_9 : out std_logic_vector( 16-1 downto 0 );
    o_10 : out std_logic_vector( 16-1 downto 0 );
    o_11 : out std_logic_vector( 16-1 downto 0 );
    o_12 : out std_logic_vector( 16-1 downto 0 );
    o_13 : out std_logic_vector( 16-1 downto 0 );
    o_14 : out std_logic_vector( 16-1 downto 0 );
    o_15 : out std_logic_vector( 16-1 downto 0 );
    o_16 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_scalar_to_vector4_x7;
architecture structural of psb3_0_scalar_to_vector4_x7 is 
  signal slice7_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 16-1 downto 0 );
  signal mux5_y_net : std_logic_vector( 256-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 16-1 downto 0 );
begin
  o_1 <= slice0_y_net;
  o_2 <= slice1_y_net;
  o_3 <= slice2_y_net;
  o_4 <= slice3_y_net;
  o_5 <= slice4_y_net;
  o_6 <= slice5_y_net;
  o_7 <= slice6_y_net;
  o_8 <= slice7_y_net;
  o_9 <= slice8_y_net;
  o_10 <= slice9_y_net;
  o_11 <= slice10_y_net;
  o_12 <= slice11_y_net;
  o_13 <= slice12_y_net;
  o_14 <= slice13_y_net;
  o_15 <= slice14_y_net;
  o_16 <= slice15_y_net;
  mux5_y_net <= i;
  slice0 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 15,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice0_y_net
  );
  slice1 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 16,
    new_msb => 31,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice1_y_net
  );
  slice2 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 32,
    new_msb => 47,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice2_y_net
  );
  slice3 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 48,
    new_msb => 63,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice3_y_net
  );
  slice4 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 64,
    new_msb => 79,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice4_y_net
  );
  slice5 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 80,
    new_msb => 95,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice5_y_net
  );
  slice6 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 96,
    new_msb => 111,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice6_y_net
  );
  slice7 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 112,
    new_msb => 127,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice7_y_net
  );
  slice8 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 128,
    new_msb => 143,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice8_y_net
  );
  slice9 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 144,
    new_msb => 159,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice9_y_net
  );
  slice10 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 160,
    new_msb => 175,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice10_y_net
  );
  slice11 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 176,
    new_msb => 191,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice11_y_net
  );
  slice12 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 192,
    new_msb => 207,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice12_y_net
  );
  slice13 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 208,
    new_msb => 223,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice13_y_net
  );
  slice14 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 224,
    new_msb => 239,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice14_y_net
  );
  slice15 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 240,
    new_msb => 255,
    x_width => 256,
    y_width => 16
  )
  port map (
    x => mux5_y_net,
    y => slice15_y_net
  );
end structural;
-- Generated from Simulink block PSB3_0/reordering extending buffer real_4/Vector Reinterpret
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_reinterpret_x10 is
  port (
    in_1 : in std_logic_vector( 16-1 downto 0 );
    in_2 : in std_logic_vector( 16-1 downto 0 );
    in_3 : in std_logic_vector( 16-1 downto 0 );
    in_4 : in std_logic_vector( 16-1 downto 0 );
    in_5 : in std_logic_vector( 16-1 downto 0 );
    in_6 : in std_logic_vector( 16-1 downto 0 );
    in_7 : in std_logic_vector( 16-1 downto 0 );
    in_8 : in std_logic_vector( 16-1 downto 0 );
    in_9 : in std_logic_vector( 16-1 downto 0 );
    in_10 : in std_logic_vector( 16-1 downto 0 );
    in_11 : in std_logic_vector( 16-1 downto 0 );
    in_12 : in std_logic_vector( 16-1 downto 0 );
    in_13 : in std_logic_vector( 16-1 downto 0 );
    in_14 : in std_logic_vector( 16-1 downto 0 );
    in_15 : in std_logic_vector( 16-1 downto 0 );
    in_16 : in std_logic_vector( 16-1 downto 0 );
    out_1 : out std_logic_vector( 16-1 downto 0 );
    out_2 : out std_logic_vector( 16-1 downto 0 );
    out_3 : out std_logic_vector( 16-1 downto 0 );
    out_4 : out std_logic_vector( 16-1 downto 0 );
    out_5 : out std_logic_vector( 16-1 downto 0 );
    out_6 : out std_logic_vector( 16-1 downto 0 );
    out_7 : out std_logic_vector( 16-1 downto 0 );
    out_8 : out std_logic_vector( 16-1 downto 0 );
    out_9 : out std_logic_vector( 16-1 downto 0 );
    out_10 : out std_logic_vector( 16-1 downto 0 );
    out_11 : out std_logic_vector( 16-1 downto 0 );
    out_12 : out std_logic_vector( 16-1 downto 0 );
    out_13 : out std_logic_vector( 16-1 downto 0 );
    out_14 : out std_logic_vector( 16-1 downto 0 );
    out_15 : out std_logic_vector( 16-1 downto 0 );
    out_16 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_vector_reinterpret_x10;
architecture structural of psb3_0_vector_reinterpret_x10 is 
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 16-1 downto 0 );
begin
  out_1 <= reinterpret0_output_port_net;
  out_2 <= reinterpret1_output_port_net;
  out_3 <= reinterpret2_output_port_net;
  out_4 <= reinterpret3_output_port_net;
  out_5 <= reinterpret4_output_port_net;
  out_6 <= reinterpret5_output_port_net;
  out_7 <= reinterpret6_output_port_net;
  out_8 <= reinterpret7_output_port_net;
  out_9 <= reinterpret8_output_port_net;
  out_10 <= reinterpret9_output_port_net;
  out_11 <= reinterpret10_output_port_net;
  out_12 <= reinterpret11_output_port_net;
  out_13 <= reinterpret12_output_port_net;
  out_14 <= reinterpret13_output_port_net;
  out_15 <= reinterpret14_output_port_net;
  out_16 <= reinterpret15_output_port_net;
  slice0_y_net <= in_1;
  slice1_y_net <= in_2;
  slice2_y_net <= in_3;
  slice3_y_net <= in_4;
  slice4_y_net <= in_5;
  slice5_y_net <= in_6;
  slice6_y_net <= in_7;
  slice7_y_net <= in_8;
  slice8_y_net <= in_9;
  slice9_y_net <= in_10;
  slice10_y_net <= in_11;
  slice11_y_net <= in_12;
  slice12_y_net <= in_13;
  slice13_y_net <= in_14;
  slice14_y_net <= in_15;
  slice15_y_net <= in_16;
  reinterpret0 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice0_y_net,
    output_port => reinterpret0_output_port_net
  );
  reinterpret1 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice1_y_net,
    output_port => reinterpret1_output_port_net
  );
  reinterpret2 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice2_y_net,
    output_port => reinterpret2_output_port_net
  );
  reinterpret3 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice3_y_net,
    output_port => reinterpret3_output_port_net
  );
  reinterpret4 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice4_y_net,
    output_port => reinterpret4_output_port_net
  );
  reinterpret5 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice5_y_net,
    output_port => reinterpret5_output_port_net
  );
  reinterpret6 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice6_y_net,
    output_port => reinterpret6_output_port_net
  );
  reinterpret7 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice7_y_net,
    output_port => reinterpret7_output_port_net
  );
  reinterpret8 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice8_y_net,
    output_port => reinterpret8_output_port_net
  );
  reinterpret9 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice9_y_net,
    output_port => reinterpret9_output_port_net
  );
  reinterpret10 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice10_y_net,
    output_port => reinterpret10_output_port_net
  );
  reinterpret11 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice11_y_net,
    output_port => reinterpret11_output_port_net
  );
  reinterpret12 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice12_y_net,
    output_port => reinterpret12_output_port_net
  );
  reinterpret13 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice13_y_net,
    output_port => reinterpret13_output_port_net
  );
  reinterpret14 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice14_y_net,
    output_port => reinterpret14_output_port_net
  );
  reinterpret15 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice15_y_net,
    output_port => reinterpret15_output_port_net
  );
end structural;
-- Generated from Simulink block PSB3_0/reordering extending buffer real_4
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_reordering_extending_buffer_real_4 is
  port (
    in_reset : in std_logic_vector( 1-1 downto 0 );
    input1 : in std_logic_vector( 16-1 downto 0 );
    input2 : in std_logic_vector( 16-1 downto 0 );
    in_tvalid : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    vec_output_1 : out std_logic_vector( 16-1 downto 0 );
    vec_output_2 : out std_logic_vector( 16-1 downto 0 );
    vec_output_3 : out std_logic_vector( 16-1 downto 0 );
    vec_output_4 : out std_logic_vector( 16-1 downto 0 );
    vec_output_5 : out std_logic_vector( 16-1 downto 0 );
    vec_output_6 : out std_logic_vector( 16-1 downto 0 );
    vec_output_7 : out std_logic_vector( 16-1 downto 0 );
    vec_output_8 : out std_logic_vector( 16-1 downto 0 );
    vec_output_9 : out std_logic_vector( 16-1 downto 0 );
    vec_output_10 : out std_logic_vector( 16-1 downto 0 );
    vec_output_11 : out std_logic_vector( 16-1 downto 0 );
    vec_output_12 : out std_logic_vector( 16-1 downto 0 );
    vec_output_13 : out std_logic_vector( 16-1 downto 0 );
    vec_output_14 : out std_logic_vector( 16-1 downto 0 );
    vec_output_15 : out std_logic_vector( 16-1 downto 0 );
    vec_output_16 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_reordering_extending_buffer_real_4;
architecture structural of psb3_0_reordering_extending_buffer_real_4 is 
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal dual_port_ram_0_doutb_net : std_logic_vector( 16-1 downto 0 );
  signal bitbasher_out_x0_net : std_logic_vector( 256-1 downto 0 );
  signal ce_net : std_logic;
  signal slice14_y_net : std_logic_vector( 16-1 downto 0 );
  signal bitbasher1_out_x0_net : std_logic_vector( 256-1 downto 0 );
  signal dual_port_ram_1_douta_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal mux7_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 16-1 downto 0 );
  signal mux3_y_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 16-1 downto 0 );
  signal dual_port_ram_0_douta_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal delay19_q_net : std_logic_vector( 1-1 downto 0 );
  signal gin_tl_reset_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal slice3_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 16-1 downto 0 );
  signal mux5_y_net : std_logic_vector( 256-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 16-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 16-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 1-1 downto 0 );
  signal single_port_ram_data_out_net : std_logic_vector( 1-1 downto 0 );
  signal delay10_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 16-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 1-1 downto 0 );
  signal constant2_op_net : std_logic_vector( 1-1 downto 0 );
  signal dual_port_ram_1_doutb_net : std_logic_vector( 16-1 downto 0 );
  signal constant_op_net : std_logic_vector( 1-1 downto 0 );
  signal we_0 : std_logic_vector( 1-1 downto 0 );
  signal delay11_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 1-1 downto 0 );
  signal addr_r_op_net : std_logic_vector( 8-1 downto 0 );
  signal delay9_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay7_q_net : std_logic_vector( 8-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 9-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 9-1 downto 0 );
  signal even_addr_w_op_net : std_logic_vector( 9-1 downto 0 );
  signal odd_addr_w_op_net : std_logic_vector( 9-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 9-1 downto 0 );
  signal mux2_y_net : std_logic_vector( 9-1 downto 0 );
  signal inverter_op_net : std_logic_vector( 1-1 downto 0 );
  signal mux4_y_net : std_logic_vector( 9-1 downto 0 );
  signal addr_control_op_net : std_logic_vector( 9-1 downto 0 );
  signal out_in_1024_out_x0_net : std_logic_vector( 9-1 downto 0 );
  signal mux3_y_net : std_logic_vector( 9-1 downto 0 );
begin
  vec_output_1 <= reinterpret0_output_port_net;
  vec_output_2 <= reinterpret1_output_port_net;
  vec_output_3 <= reinterpret2_output_port_net;
  vec_output_4 <= reinterpret3_output_port_net;
  vec_output_5 <= reinterpret4_output_port_net;
  vec_output_6 <= reinterpret5_output_port_net;
  vec_output_7 <= reinterpret6_output_port_net;
  vec_output_8 <= reinterpret7_output_port_net;
  vec_output_9 <= reinterpret8_output_port_net;
  vec_output_10 <= reinterpret9_output_port_net;
  vec_output_11 <= reinterpret10_output_port_net;
  vec_output_12 <= reinterpret11_output_port_net;
  vec_output_13 <= reinterpret12_output_port_net;
  vec_output_14 <= reinterpret13_output_port_net;
  vec_output_15 <= reinterpret14_output_port_net;
  vec_output_16 <= reinterpret15_output_port_net;
  gin_tl_reset_net <= in_reset;
  mux3_y_net_x0 <= input1;
  mux7_y_net <= input2;
  delay19_q_net <= in_tvalid;
  clk_net <= clk_1;
  ce_net <= ce_1;
  scalar_to_vector4 : entity xil_defaultlib.psb3_0_scalar_to_vector4_x7 
  port map (
    i => mux5_y_net,
    o_1 => slice0_y_net,
    o_2 => slice1_y_net,
    o_3 => slice2_y_net,
    o_4 => slice3_y_net,
    o_5 => slice4_y_net,
    o_6 => slice5_y_net,
    o_7 => slice6_y_net,
    o_8 => slice7_y_net,
    o_9 => slice8_y_net,
    o_10 => slice9_y_net,
    o_11 => slice10_y_net,
    o_12 => slice11_y_net,
    o_13 => slice12_y_net,
    o_14 => slice13_y_net,
    o_15 => slice14_y_net,
    o_16 => slice15_y_net
  );
  vector_reinterpret : entity xil_defaultlib.psb3_0_vector_reinterpret_x10 
  port map (
    in_1 => slice0_y_net,
    in_2 => slice1_y_net,
    in_3 => slice2_y_net,
    in_4 => slice3_y_net,
    in_5 => slice4_y_net,
    in_6 => slice5_y_net,
    in_7 => slice6_y_net,
    in_8 => slice7_y_net,
    in_9 => slice8_y_net,
    in_10 => slice9_y_net,
    in_11 => slice10_y_net,
    in_12 => slice11_y_net,
    in_13 => slice12_y_net,
    in_14 => slice13_y_net,
    in_15 => slice14_y_net,
    in_16 => slice15_y_net,
    out_1 => reinterpret0_output_port_net,
    out_2 => reinterpret1_output_port_net,
    out_3 => reinterpret2_output_port_net,
    out_4 => reinterpret3_output_port_net,
    out_5 => reinterpret4_output_port_net,
    out_6 => reinterpret5_output_port_net,
    out_7 => reinterpret6_output_port_net,
    out_8 => reinterpret7_output_port_net,
    out_9 => reinterpret8_output_port_net,
    out_10 => reinterpret9_output_port_net,
    out_11 => reinterpret10_output_port_net,
    out_12 => reinterpret11_output_port_net,
    out_13 => reinterpret12_output_port_net,
    out_14 => reinterpret13_output_port_net,
    out_15 => reinterpret14_output_port_net,
    out_16 => reinterpret15_output_port_net
  );
  bitbasher : entity xil_defaultlib.sysgen_bitbasher_4648460ba6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    a => dual_port_ram_0_douta_net,
    b => dual_port_ram_0_doutb_net,
    out_x0 => bitbasher_out_x0_net
  );
  bitbasher1 : entity xil_defaultlib.sysgen_bitbasher_4648460ba6 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    a => dual_port_ram_1_douta_net,
    b => dual_port_ram_1_doutb_net,
    out_x0 => bitbasher1_out_x0_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_de9059c03f 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_71e89d757c 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  constant2 : entity xil_defaultlib.sysgen_constant_71e89d757c 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant2_op_net
  );
  delay : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => single_port_ram_data_out_net,
    clk => clk_net,
    ce => ce_net,
    q => we_0
  );
  delay1 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 16
  )
  port map (
    en => '1',
    rst => '0',
    d => mux3_y_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay10 : entity xil_defaultlib.sysgen_delay_906db00812 
  port map (
    clr => '0',
    d => constant1_op_net,
    rst => gin_tl_reset_net,
    clk => clk_net,
    ce => ce_net,
    q => delay10_q_net
  );
  delay11 : entity xil_defaultlib.sysgen_delay_906db00812 
  port map (
    clr => '0',
    d => constant2_op_net,
    rst => gin_tl_reset_net,
    clk => clk_net,
    ce => ce_net,
    q => delay11_q_net
  );
  delay2 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 16
  )
  port map (
    en => '1',
    rst => '0',
    d => mux7_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay3 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => we_0,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  delay4 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => inverter_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net
  );
  delay5 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 9
  )
  port map (
    en => '1',
    rst => '0',
    d => even_addr_w_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  delay6 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 9
  )
  port map (
    en => '1',
    rst => '0',
    d => odd_addr_w_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay6_q_net
  );
  delay7 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 8
  )
  port map (
    en => '1',
    rst => '0',
    d => addr_r_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay7_q_net
  );
  delay9 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay9_q_net
  );
  dual_port_ram_0 : entity xil_defaultlib.psb3_0_xltdpram 
  generic map (
    addr_width_b => 9,
    clocking_mode => "common_clock",
    data_width_b => 16,
    latency => 1,
    mem_init_file => "xpm_c5fd30_vivado.mem",
    mem_size => 8192,
    mem_type => "block",
    read_reset_a => "0",
    read_reset_b => "0",
    width => 16,
    width_addr => 9,
    write_mode_a => "read_first",
    write_mode_b => "read_first"
  )
  port map (
    ena => "1",
    rsta => "0",
    rstb => "0",
    addra => mux1_y_net,
    dina => delay1_q_net,
    wea => delay3_q_net,
    addrb => mux2_y_net,
    dinb => delay2_q_net,
    web => delay3_q_net,
    enb => delay11_q_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dual_port_ram_0_douta_net,
    doutb => dual_port_ram_0_doutb_net
  );
  dual_port_ram_1 : entity xil_defaultlib.psb3_0_xltdpram 
  generic map (
    addr_width_b => 9,
    clocking_mode => "common_clock",
    data_width_b => 16,
    latency => 1,
    mem_init_file => "xpm_c5fd30_vivado.mem",
    mem_size => 8192,
    mem_type => "block",
    read_reset_a => "0",
    read_reset_b => "0",
    width => 16,
    width_addr => 9,
    write_mode_a => "read_first",
    write_mode_b => "read_first"
  )
  port map (
    ena => "1",
    rsta => "0",
    rstb => "0",
    addra => mux3_y_net,
    dina => delay1_q_net,
    wea => delay4_q_net,
    addrb => mux4_y_net,
    dinb => delay2_q_net,
    web => delay4_q_net,
    enb => delay10_q_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dual_port_ram_1_douta_net,
    doutb => dual_port_ram_1_doutb_net
  );
  inverter : entity xil_defaultlib.sysgen_inverter_ac5174c184 
  port map (
    clr => '0',
    ip => single_port_ram_data_out_net,
    clk => clk_net,
    ce => ce_net,
    op => inverter_op_net
  );
  mux1 : entity xil_defaultlib.sysgen_mux_303302b1e4 
  port map (
    clr => '0',
    sel => we_0,
    d0 => delay7_q_net,
    d1 => delay5_q_net,
    clk => clk_net,
    ce => ce_net,
    y => mux1_y_net
  );
  mux2 : entity xil_defaultlib.sysgen_mux_c7d0cfa098 
  port map (
    clr => '0',
    sel => we_0,
    d0 => out_in_1024_out_x0_net,
    d1 => delay6_q_net,
    clk => clk_net,
    ce => ce_net,
    y => mux2_y_net
  );
  mux3 : entity xil_defaultlib.sysgen_mux_303302b1e4 
  port map (
    clr => '0',
    sel => inverter_op_net,
    d0 => delay7_q_net,
    d1 => delay5_q_net,
    clk => clk_net,
    ce => ce_net,
    y => mux3_y_net
  );
  mux4 : entity xil_defaultlib.sysgen_mux_c7d0cfa098 
  port map (
    clr => '0',
    sel => inverter_op_net,
    d0 => out_in_1024_out_x0_net,
    d1 => delay6_q_net,
    clk => clk_net,
    ce => ce_net,
    y => mux4_y_net
  );
  mux5 : entity xil_defaultlib.sysgen_mux_1f606cf16b 
  port map (
    clr => '0',
    sel => delay9_q_net,
    d0 => bitbasher_out_x0_net,
    d1 => bitbasher1_out_x0_net,
    clk => clk_net,
    ce => ce_net,
    y => mux5_y_net
  );
  single_port_ram : entity xil_defaultlib.psb3_0_xlspram 
  generic map (
    init_value => b"0",
    latency => 1,
    mem_init_file => "xpm_95b604_vivado.mem",
    mem_size => 512,
    mem_type => "block",
    read_reset_val => "0",
    width => 1,
    width_addr => 9,
    write_mode_a => "read_first",
    xpm_lat => 1
  )
  port map (
    en => "1",
    rst => "0",
    addr => addr_control_op_net,
    data_in => constant_op_net,
    we => constant_op_net,
    clk => clk_net,
    ce => ce_net,
    data_out => single_port_ram_data_out_net
  );
  addr_control : entity xil_defaultlib.psb3_0_xlcounter_free 
  generic map (
    core_name0 => "psb3_0_c_counter_binary_v12_0_i4",
    op_arith => xlUnsigned,
    op_width => 9
  )
  port map (
    clr => '0',
    rst => gin_tl_reset_net,
    en => delay19_q_net,
    clk => clk_net,
    ce => ce_net,
    op => addr_control_op_net
  );
  addr_r : entity xil_defaultlib.psb3_0_xlcounter_free 
  generic map (
    core_name0 => "psb3_0_c_counter_binary_v12_0_i3",
    op_arith => xlUnsigned,
    op_width => 8
  )
  port map (
    clr => '0',
    rst => gin_tl_reset_net,
    en => delay19_q_net,
    clk => clk_net,
    ce => ce_net,
    op => addr_r_op_net
  );
  even_addr_w : entity xil_defaultlib.psb3_0_xlcounter_free 
  generic map (
    core_name0 => "psb3_0_c_counter_binary_v12_0_i5",
    op_arith => xlUnsigned,
    op_width => 9
  )
  port map (
    clr => '0',
    rst => gin_tl_reset_net,
    en => delay19_q_net,
    clk => clk_net,
    ce => ce_net,
    op => even_addr_w_op_net
  );
  odd_addr_w : entity xil_defaultlib.psb3_0_xlcounter_free 
  generic map (
    core_name0 => "psb3_0_c_counter_binary_v12_0_i6",
    op_arith => xlUnsigned,
    op_width => 9
  )
  port map (
    clr => '0',
    rst => gin_tl_reset_net,
    en => delay19_q_net,
    clk => clk_net,
    ce => ce_net,
    op => odd_addr_w_op_net
  );
  out_in_1024 : entity xil_defaultlib.sysgen_bitbasher_a62d2ce679 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in_x0 => delay7_q_net,
    out_x0 => out_in_1024_out_x0_net
  );
end structural;
-- Generated from Simulink block PSB3_0/vector IFFT/Vector FFT
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_fft is
  port (
    i_re_1 : in std_logic_vector( 17-1 downto 0 );
    i_im_1 : in std_logic_vector( 17-1 downto 0 );
    vi : in std_logic_vector( 1-1 downto 0 );
    si : in std_logic_vector( 11-1 downto 0 );
    i_re_2 : in std_logic_vector( 17-1 downto 0 );
    i_re_3 : in std_logic_vector( 17-1 downto 0 );
    i_re_4 : in std_logic_vector( 17-1 downto 0 );
    i_re_5 : in std_logic_vector( 17-1 downto 0 );
    i_re_6 : in std_logic_vector( 17-1 downto 0 );
    i_re_7 : in std_logic_vector( 17-1 downto 0 );
    i_re_8 : in std_logic_vector( 17-1 downto 0 );
    i_im_2 : in std_logic_vector( 17-1 downto 0 );
    i_im_3 : in std_logic_vector( 17-1 downto 0 );
    i_im_4 : in std_logic_vector( 17-1 downto 0 );
    i_im_5 : in std_logic_vector( 17-1 downto 0 );
    i_im_6 : in std_logic_vector( 17-1 downto 0 );
    i_im_7 : in std_logic_vector( 17-1 downto 0 );
    i_im_8 : in std_logic_vector( 17-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    o_re_1 : out std_logic_vector( 20-1 downto 0 );
    o_im_1 : out std_logic_vector( 20-1 downto 0 );
    vo : out std_logic;
    o_re_2 : out std_logic_vector( 20-1 downto 0 );
    o_re_3 : out std_logic_vector( 20-1 downto 0 );
    o_re_4 : out std_logic_vector( 20-1 downto 0 );
    o_re_5 : out std_logic_vector( 20-1 downto 0 );
    o_re_6 : out std_logic_vector( 20-1 downto 0 );
    o_re_7 : out std_logic_vector( 20-1 downto 0 );
    o_re_8 : out std_logic_vector( 20-1 downto 0 );
    o_im_2 : out std_logic_vector( 20-1 downto 0 );
    o_im_3 : out std_logic_vector( 20-1 downto 0 );
    o_im_4 : out std_logic_vector( 20-1 downto 0 );
    o_im_5 : out std_logic_vector( 20-1 downto 0 );
    o_im_6 : out std_logic_vector( 20-1 downto 0 );
    o_im_7 : out std_logic_vector( 20-1 downto 0 );
    o_im_8 : out std_logic_vector( 20-1 downto 0 )
  );
end psb3_0_vector_fft;
architecture structural of psb3_0_vector_fft is 
  signal reinterpret25_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal mux2_y_net : std_logic_vector( 17-1 downto 0 );
  signal reinterpret19_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal reinterpret17_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal delay11_q_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret31_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal reinterpret20_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal reinterpret30_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal test_systolicfft_vhdl_black_box_vo_net : std_logic;
  signal constant15_op_net : std_logic_vector( 11-1 downto 0 );
  signal reinterpret18_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal reinterpret23_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal reinterpret24_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal reinterpret26_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal reinterpret21_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal reinterpret27_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal reinterpret29_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal reinterpret22_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal reinterpret16_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal reinterpret28_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal mux27_y_net : std_logic_vector( 17-1 downto 0 );
  signal mux33_y_net : std_logic_vector( 17-1 downto 0 );
  signal mux45_y_net : std_logic_vector( 17-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 11-1 downto 0 );
  signal mux54_y_net : std_logic_vector( 17-1 downto 0 );
  signal ce_net : std_logic;
  signal reinterpret1_output_port_net : std_logic_vector( 17-1 downto 0 );
  signal mux53_y_net : std_logic_vector( 17-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 17-1 downto 0 );
  signal mux46_y_net : std_logic_vector( 17-1 downto 0 );
  signal reinterpret0_output_port_net : std_logic_vector( 17-1 downto 0 );
  signal mux42_y_net : std_logic_vector( 17-1 downto 0 );
  signal mux38_y_net : std_logic_vector( 17-1 downto 0 );
  signal mux30_y_net : std_logic_vector( 17-1 downto 0 );
  signal mux37_y_net : std_logic_vector( 17-1 downto 0 );
  signal mux41_y_net : std_logic_vector( 17-1 downto 0 );
  signal mux49_y_net : std_logic_vector( 17-1 downto 0 );
  signal mux34_y_net : std_logic_vector( 17-1 downto 0 );
  signal clk_net : std_logic;
  signal delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux50_y_net : std_logic_vector( 17-1 downto 0 );
  signal mux29_y_net : std_logic_vector( 17-1 downto 0 );
  signal concat8_y_net : std_logic_vector( 272-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 17-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 17-1 downto 0 );
  signal reinterpret10_output_port_net : std_logic_vector( 17-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 17-1 downto 0 );
  signal reinterpret6_output_port_net : std_logic_vector( 17-1 downto 0 );
  signal test_systolicfft_vhdl_black_box_so_net : std_logic_vector( 11-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 17-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 17-1 downto 0 );
  signal test_systolicfft_vhdl_black_box_o_net : std_logic_vector( 320-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 17-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 17-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 17-1 downto 0 );
  signal concat4_y_net : std_logic_vector( 34-1 downto 0 );
  signal reinterpret12_output_port_net : std_logic_vector( 17-1 downto 0 );
  signal concat2_y_net : std_logic_vector( 34-1 downto 0 );
  signal concat0_y_net : std_logic_vector( 34-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 17-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 17-1 downto 0 );
  signal concat1_y_net : std_logic_vector( 34-1 downto 0 );
  signal concat3_y_net : std_logic_vector( 34-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 34-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 34-1 downto 0 );
  signal concat5_y_net : std_logic_vector( 34-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 34-1 downto 0 );
  signal concat6_y_net : std_logic_vector( 34-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 34-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 34-1 downto 0 );
  signal concat7_y_net : std_logic_vector( 34-1 downto 0 );
  signal delay7_q_net : std_logic_vector( 34-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 40-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 20-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 40-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 20-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 20-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 20-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 40-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 20-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 40-1 downto 0 );
  signal delay9_q_net : std_logic_vector( 34-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 34-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 40-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 40-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 40-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 40-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 20-1 downto 0 );
  signal slice23_y_net : std_logic_vector( 20-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 20-1 downto 0 );
  signal slice22_y_net : std_logic_vector( 20-1 downto 0 );
  signal slice20_y_net : std_logic_vector( 20-1 downto 0 );
  signal slice19_y_net : std_logic_vector( 20-1 downto 0 );
  signal slice18_y_net : std_logic_vector( 20-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 20-1 downto 0 );
  signal slice17_y_net : std_logic_vector( 20-1 downto 0 );
  signal slice16_y_net : std_logic_vector( 20-1 downto 0 );
  signal slice21_y_net : std_logic_vector( 20-1 downto 0 );
begin
  o_re_1 <= reinterpret16_output_port_net;
  o_im_1 <= reinterpret24_output_port_net;
  vo <= test_systolicfft_vhdl_black_box_vo_net;
  o_re_2 <= reinterpret17_output_port_net;
  o_re_3 <= reinterpret18_output_port_net;
  o_re_4 <= reinterpret19_output_port_net;
  o_re_5 <= reinterpret20_output_port_net;
  o_re_6 <= reinterpret21_output_port_net;
  o_re_7 <= reinterpret22_output_port_net;
  o_re_8 <= reinterpret23_output_port_net;
  o_im_2 <= reinterpret25_output_port_net;
  o_im_3 <= reinterpret26_output_port_net;
  o_im_4 <= reinterpret27_output_port_net;
  o_im_5 <= reinterpret28_output_port_net;
  o_im_6 <= reinterpret29_output_port_net;
  o_im_7 <= reinterpret30_output_port_net;
  o_im_8 <= reinterpret31_output_port_net;
  mux27_y_net <= i_re_1;
  mux2_y_net <= i_im_1;
  delay11_q_net <= vi;
  constant15_op_net <= si;
  mux30_y_net <= i_re_2;
  mux34_y_net <= i_re_3;
  mux38_y_net <= i_re_4;
  mux42_y_net <= i_re_5;
  mux46_y_net <= i_re_6;
  mux50_y_net <= i_re_7;
  mux54_y_net <= i_re_8;
  mux29_y_net <= i_im_2;
  mux33_y_net <= i_im_3;
  mux37_y_net <= i_im_4;
  mux41_y_net <= i_im_5;
  mux45_y_net <= i_im_6;
  mux49_y_net <= i_im_7;
  mux53_y_net <= i_im_8;
  clk_net <= clk_1;
  ce_net <= ce_1;
  delay : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 4,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay11_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_q_net
  );
  delay1 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 4,
    reg_retiming => 0,
    reset => 0,
    width => 11
  )
  port map (
    en => '1',
    rst => '0',
    d => constant15_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  reinterpret0 : entity xil_defaultlib.sysgen_reinterpret_432d320890 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => mux2_y_net,
    output_port => reinterpret0_output_port_net
  );
  reinterpret1 : entity xil_defaultlib.sysgen_reinterpret_432d320890 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => mux29_y_net,
    output_port => reinterpret1_output_port_net
  );
  reinterpret2 : entity xil_defaultlib.sysgen_reinterpret_432d320890 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => mux33_y_net,
    output_port => reinterpret2_output_port_net
  );
  test_systolicfft_vhdl_black_box : entity xil_defaultlib.WRAPPER_VECTOR_FFT_b8a7010354694656355591d9cada5b52 
  generic map (
    BRAM_THRESHOLD => 258,
    DSP48E => 2,
    I_high => 1,
    I_low => -15,
    L2N => 11,
    N => 2048,
    O_high => 4,
    O_low => -15,
    SSR => 8,
    W_high => 1,
    W_low => -17
  )
  port map (
    i => concat8_y_net,
    vi => delay_q_net(0),
    si => delay1_q_net,
    CLK => clk_net,
    CE => ce_net,
    o => test_systolicfft_vhdl_black_box_o_net,
    vo => test_systolicfft_vhdl_black_box_vo_net,
    so => test_systolicfft_vhdl_black_box_so_net
  );
  reinterpret3 : entity xil_defaultlib.sysgen_reinterpret_432d320890 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => mux37_y_net,
    output_port => reinterpret3_output_port_net
  );
  reinterpret4 : entity xil_defaultlib.sysgen_reinterpret_432d320890 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => mux41_y_net,
    output_port => reinterpret4_output_port_net
  );
  reinterpret5 : entity xil_defaultlib.sysgen_reinterpret_432d320890 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => mux45_y_net,
    output_port => reinterpret5_output_port_net
  );
  reinterpret6 : entity xil_defaultlib.sysgen_reinterpret_432d320890 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => mux49_y_net,
    output_port => reinterpret6_output_port_net
  );
  reinterpret7 : entity xil_defaultlib.sysgen_reinterpret_432d320890 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => mux53_y_net,
    output_port => reinterpret7_output_port_net
  );
  reinterpret8 : entity xil_defaultlib.sysgen_reinterpret_432d320890 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => mux27_y_net,
    output_port => reinterpret8_output_port_net
  );
  reinterpret9 : entity xil_defaultlib.sysgen_reinterpret_432d320890 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => mux30_y_net,
    output_port => reinterpret9_output_port_net
  );
  reinterpret10 : entity xil_defaultlib.sysgen_reinterpret_432d320890 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => mux34_y_net,
    output_port => reinterpret10_output_port_net
  );
  reinterpret11 : entity xil_defaultlib.sysgen_reinterpret_432d320890 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => mux38_y_net,
    output_port => reinterpret11_output_port_net
  );
  reinterpret12 : entity xil_defaultlib.sysgen_reinterpret_432d320890 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => mux42_y_net,
    output_port => reinterpret12_output_port_net
  );
  reinterpret13 : entity xil_defaultlib.sysgen_reinterpret_432d320890 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => mux46_y_net,
    output_port => reinterpret13_output_port_net
  );
  reinterpret14 : entity xil_defaultlib.sysgen_reinterpret_432d320890 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => mux50_y_net,
    output_port => reinterpret14_output_port_net
  );
  reinterpret15 : entity xil_defaultlib.sysgen_reinterpret_432d320890 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => mux54_y_net,
    output_port => reinterpret15_output_port_net
  );
  concat0 : entity xil_defaultlib.sysgen_concat_1b398cb1a1 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => reinterpret0_output_port_net,
    in1 => reinterpret8_output_port_net,
    y => concat0_y_net
  );
  concat1 : entity xil_defaultlib.sysgen_concat_1b398cb1a1 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => reinterpret1_output_port_net,
    in1 => reinterpret9_output_port_net,
    y => concat1_y_net
  );
  concat2 : entity xil_defaultlib.sysgen_concat_1b398cb1a1 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => reinterpret2_output_port_net,
    in1 => reinterpret10_output_port_net,
    y => concat2_y_net
  );
  concat3 : entity xil_defaultlib.sysgen_concat_1b398cb1a1 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => reinterpret3_output_port_net,
    in1 => reinterpret11_output_port_net,
    y => concat3_y_net
  );
  concat4 : entity xil_defaultlib.sysgen_concat_1b398cb1a1 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => reinterpret4_output_port_net,
    in1 => reinterpret12_output_port_net,
    y => concat4_y_net
  );
  concat5 : entity xil_defaultlib.sysgen_concat_1b398cb1a1 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => reinterpret5_output_port_net,
    in1 => reinterpret13_output_port_net,
    y => concat5_y_net
  );
  concat6 : entity xil_defaultlib.sysgen_concat_1b398cb1a1 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => reinterpret6_output_port_net,
    in1 => reinterpret14_output_port_net,
    y => concat6_y_net
  );
  concat7 : entity xil_defaultlib.sysgen_concat_1b398cb1a1 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => reinterpret7_output_port_net,
    in1 => reinterpret15_output_port_net,
    y => concat7_y_net
  );
  delay2 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 4,
    reg_retiming => 0,
    reset => 0,
    width => 34
  )
  port map (
    en => '1',
    rst => '0',
    d => concat0_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay3 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 4,
    reg_retiming => 0,
    reset => 0,
    width => 34
  )
  port map (
    en => '1',
    rst => '0',
    d => concat1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  delay4 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 4,
    reg_retiming => 0,
    reset => 0,
    width => 34
  )
  port map (
    en => '1',
    rst => '0',
    d => concat2_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net
  );
  delay5 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 4,
    reg_retiming => 0,
    reset => 0,
    width => 34
  )
  port map (
    en => '1',
    rst => '0',
    d => concat3_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  delay6 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 4,
    reg_retiming => 0,
    reset => 0,
    width => 34
  )
  port map (
    en => '1',
    rst => '0',
    d => concat4_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay6_q_net
  );
  delay7 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 4,
    reg_retiming => 0,
    reset => 0,
    width => 34
  )
  port map (
    en => '1',
    rst => '0',
    d => concat5_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay7_q_net
  );
  delay8 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 4,
    reg_retiming => 0,
    reset => 0,
    width => 34
  )
  port map (
    en => '1',
    rst => '0',
    d => concat6_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay8_q_net
  );
  delay9 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 4,
    reg_retiming => 0,
    reset => 0,
    width => 34
  )
  port map (
    en => '1',
    rst => '0',
    d => concat7_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay9_q_net
  );
  concat8 : entity xil_defaultlib.sysgen_concat_546535937a 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => delay9_q_net,
    in1 => delay8_q_net,
    in2 => delay7_q_net,
    in3 => delay6_q_net,
    in4 => delay5_q_net,
    in5 => delay4_q_net,
    in6 => delay3_q_net,
    in7 => delay2_q_net,
    y => concat8_y_net
  );
  slice0 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 39,
    x_width => 320,
    y_width => 40
  )
  port map (
    x => test_systolicfft_vhdl_black_box_o_net,
    y => slice0_y_net
  );
  slice1 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 40,
    new_msb => 79,
    x_width => 320,
    y_width => 40
  )
  port map (
    x => test_systolicfft_vhdl_black_box_o_net,
    y => slice1_y_net
  );
  slice2 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 80,
    new_msb => 119,
    x_width => 320,
    y_width => 40
  )
  port map (
    x => test_systolicfft_vhdl_black_box_o_net,
    y => slice2_y_net
  );
  slice3 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 120,
    new_msb => 159,
    x_width => 320,
    y_width => 40
  )
  port map (
    x => test_systolicfft_vhdl_black_box_o_net,
    y => slice3_y_net
  );
  slice4 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 160,
    new_msb => 199,
    x_width => 320,
    y_width => 40
  )
  port map (
    x => test_systolicfft_vhdl_black_box_o_net,
    y => slice4_y_net
  );
  slice5 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 200,
    new_msb => 239,
    x_width => 320,
    y_width => 40
  )
  port map (
    x => test_systolicfft_vhdl_black_box_o_net,
    y => slice5_y_net
  );
  slice6 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 240,
    new_msb => 279,
    x_width => 320,
    y_width => 40
  )
  port map (
    x => test_systolicfft_vhdl_black_box_o_net,
    y => slice6_y_net
  );
  slice7 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 280,
    new_msb => 319,
    x_width => 320,
    y_width => 40
  )
  port map (
    x => test_systolicfft_vhdl_black_box_o_net,
    y => slice7_y_net
  );
  slice8 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 19,
    x_width => 40,
    y_width => 20
  )
  port map (
    x => slice0_y_net,
    y => slice8_y_net
  );
  slice9 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 19,
    x_width => 40,
    y_width => 20
  )
  port map (
    x => slice1_y_net,
    y => slice9_y_net
  );
  slice10 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 19,
    x_width => 40,
    y_width => 20
  )
  port map (
    x => slice2_y_net,
    y => slice10_y_net
  );
  slice11 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 19,
    x_width => 40,
    y_width => 20
  )
  port map (
    x => slice3_y_net,
    y => slice11_y_net
  );
  slice12 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 19,
    x_width => 40,
    y_width => 20
  )
  port map (
    x => slice4_y_net,
    y => slice12_y_net
  );
  slice13 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 19,
    x_width => 40,
    y_width => 20
  )
  port map (
    x => slice5_y_net,
    y => slice13_y_net
  );
  slice14 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 19,
    x_width => 40,
    y_width => 20
  )
  port map (
    x => slice6_y_net,
    y => slice14_y_net
  );
  slice15 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 0,
    new_msb => 19,
    x_width => 40,
    y_width => 20
  )
  port map (
    x => slice7_y_net,
    y => slice15_y_net
  );
  slice16 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 20,
    new_msb => 39,
    x_width => 40,
    y_width => 20
  )
  port map (
    x => slice0_y_net,
    y => slice16_y_net
  );
  slice17 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 20,
    new_msb => 39,
    x_width => 40,
    y_width => 20
  )
  port map (
    x => slice1_y_net,
    y => slice17_y_net
  );
  slice18 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 20,
    new_msb => 39,
    x_width => 40,
    y_width => 20
  )
  port map (
    x => slice2_y_net,
    y => slice18_y_net
  );
  slice19 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 20,
    new_msb => 39,
    x_width => 40,
    y_width => 20
  )
  port map (
    x => slice3_y_net,
    y => slice19_y_net
  );
  slice20 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 20,
    new_msb => 39,
    x_width => 40,
    y_width => 20
  )
  port map (
    x => slice4_y_net,
    y => slice20_y_net
  );
  slice21 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 20,
    new_msb => 39,
    x_width => 40,
    y_width => 20
  )
  port map (
    x => slice5_y_net,
    y => slice21_y_net
  );
  slice22 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 20,
    new_msb => 39,
    x_width => 40,
    y_width => 20
  )
  port map (
    x => slice6_y_net,
    y => slice22_y_net
  );
  slice23 : entity xil_defaultlib.psb3_0_xlslice 
  generic map (
    new_lsb => 20,
    new_msb => 39,
    x_width => 40,
    y_width => 20
  )
  port map (
    x => slice7_y_net,
    y => slice23_y_net
  );
  reinterpret16 : entity xil_defaultlib.sysgen_reinterpret_bcba3ccfb1 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice8_y_net,
    output_port => reinterpret16_output_port_net
  );
  reinterpret17 : entity xil_defaultlib.sysgen_reinterpret_bcba3ccfb1 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice9_y_net,
    output_port => reinterpret17_output_port_net
  );
  reinterpret18 : entity xil_defaultlib.sysgen_reinterpret_bcba3ccfb1 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice10_y_net,
    output_port => reinterpret18_output_port_net
  );
  reinterpret19 : entity xil_defaultlib.sysgen_reinterpret_bcba3ccfb1 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice11_y_net,
    output_port => reinterpret19_output_port_net
  );
  reinterpret20 : entity xil_defaultlib.sysgen_reinterpret_bcba3ccfb1 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice12_y_net,
    output_port => reinterpret20_output_port_net
  );
  reinterpret21 : entity xil_defaultlib.sysgen_reinterpret_bcba3ccfb1 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice13_y_net,
    output_port => reinterpret21_output_port_net
  );
  reinterpret22 : entity xil_defaultlib.sysgen_reinterpret_bcba3ccfb1 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice14_y_net,
    output_port => reinterpret22_output_port_net
  );
  reinterpret23 : entity xil_defaultlib.sysgen_reinterpret_bcba3ccfb1 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice15_y_net,
    output_port => reinterpret23_output_port_net
  );
  reinterpret24 : entity xil_defaultlib.sysgen_reinterpret_bcba3ccfb1 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice16_y_net,
    output_port => reinterpret24_output_port_net
  );
  reinterpret25 : entity xil_defaultlib.sysgen_reinterpret_bcba3ccfb1 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice17_y_net,
    output_port => reinterpret25_output_port_net
  );
  reinterpret26 : entity xil_defaultlib.sysgen_reinterpret_bcba3ccfb1 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice18_y_net,
    output_port => reinterpret26_output_port_net
  );
  reinterpret27 : entity xil_defaultlib.sysgen_reinterpret_bcba3ccfb1 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice19_y_net,
    output_port => reinterpret27_output_port_net
  );
  reinterpret28 : entity xil_defaultlib.sysgen_reinterpret_bcba3ccfb1 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice20_y_net,
    output_port => reinterpret28_output_port_net
  );
  reinterpret29 : entity xil_defaultlib.sysgen_reinterpret_bcba3ccfb1 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice21_y_net,
    output_port => reinterpret29_output_port_net
  );
  reinterpret30 : entity xil_defaultlib.sysgen_reinterpret_bcba3ccfb1 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice22_y_net,
    output_port => reinterpret30_output_port_net
  );
  reinterpret31 : entity xil_defaultlib.sysgen_reinterpret_bcba3ccfb1 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice23_y_net,
    output_port => reinterpret31_output_port_net
  );
end structural;
-- Generated from Simulink block PSB3_0/vector IFFT
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_vector_ifft is
  port (
    i_re_1 : in std_logic_vector( 17-1 downto 0 );
    i_im_1 : in std_logic_vector( 17-1 downto 0 );
    vi : in std_logic_vector( 1-1 downto 0 );
    si : in std_logic_vector( 11-1 downto 0 );
    i_re_2 : in std_logic_vector( 17-1 downto 0 );
    i_re_3 : in std_logic_vector( 17-1 downto 0 );
    i_re_4 : in std_logic_vector( 17-1 downto 0 );
    i_re_5 : in std_logic_vector( 17-1 downto 0 );
    i_re_6 : in std_logic_vector( 17-1 downto 0 );
    i_re_7 : in std_logic_vector( 17-1 downto 0 );
    i_re_8 : in std_logic_vector( 17-1 downto 0 );
    i_im_2 : in std_logic_vector( 17-1 downto 0 );
    i_im_3 : in std_logic_vector( 17-1 downto 0 );
    i_im_4 : in std_logic_vector( 17-1 downto 0 );
    i_im_5 : in std_logic_vector( 17-1 downto 0 );
    i_im_6 : in std_logic_vector( 17-1 downto 0 );
    i_im_7 : in std_logic_vector( 17-1 downto 0 );
    i_im_8 : in std_logic_vector( 17-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    o_re_1 : out std_logic_vector( 20-1 downto 0 );
    o_im_1 : out std_logic_vector( 20-1 downto 0 );
    vo : out std_logic;
    o_re_2 : out std_logic_vector( 20-1 downto 0 );
    o_re_3 : out std_logic_vector( 20-1 downto 0 );
    o_re_4 : out std_logic_vector( 20-1 downto 0 );
    o_re_5 : out std_logic_vector( 20-1 downto 0 );
    o_re_6 : out std_logic_vector( 20-1 downto 0 );
    o_re_7 : out std_logic_vector( 20-1 downto 0 );
    o_re_8 : out std_logic_vector( 20-1 downto 0 );
    o_im_2 : out std_logic_vector( 20-1 downto 0 );
    o_im_3 : out std_logic_vector( 20-1 downto 0 );
    o_im_4 : out std_logic_vector( 20-1 downto 0 );
    o_im_5 : out std_logic_vector( 20-1 downto 0 );
    o_im_6 : out std_logic_vector( 20-1 downto 0 );
    o_im_7 : out std_logic_vector( 20-1 downto 0 );
    o_im_8 : out std_logic_vector( 20-1 downto 0 )
  );
end psb3_0_vector_ifft;
architecture structural of psb3_0_vector_ifft is 
  signal reinterpret24_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal reinterpret16_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal reinterpret25_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal reinterpret26_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal reinterpret27_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal reinterpret30_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal reinterpret29_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal test_systolicfft_vhdl_black_box_vo_net : std_logic;
  signal reinterpret28_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal reinterpret21_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal reinterpret18_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal reinterpret17_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal reinterpret22_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal mux27_y_net : std_logic_vector( 17-1 downto 0 );
  signal constant15_op_net : std_logic_vector( 11-1 downto 0 );
  signal clk_net : std_logic;
  signal mux29_y_net : std_logic_vector( 17-1 downto 0 );
  signal mux41_y_net : std_logic_vector( 17-1 downto 0 );
  signal reinterpret19_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal mux33_y_net : std_logic_vector( 17-1 downto 0 );
  signal reinterpret23_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal mux53_y_net : std_logic_vector( 17-1 downto 0 );
  signal mux42_y_net : std_logic_vector( 17-1 downto 0 );
  signal mux38_y_net : std_logic_vector( 17-1 downto 0 );
  signal mux54_y_net : std_logic_vector( 17-1 downto 0 );
  signal ce_net : std_logic;
  signal reinterpret20_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal mux37_y_net : std_logic_vector( 17-1 downto 0 );
  signal mux49_y_net : std_logic_vector( 17-1 downto 0 );
  signal mux2_y_net : std_logic_vector( 17-1 downto 0 );
  signal mux30_y_net : std_logic_vector( 17-1 downto 0 );
  signal mux34_y_net : std_logic_vector( 17-1 downto 0 );
  signal reinterpret31_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal mux50_y_net : std_logic_vector( 17-1 downto 0 );
  signal mux46_y_net : std_logic_vector( 17-1 downto 0 );
  signal delay11_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux45_y_net : std_logic_vector( 17-1 downto 0 );
begin
  o_re_1 <= reinterpret24_output_port_net;
  o_im_1 <= reinterpret16_output_port_net;
  vo <= test_systolicfft_vhdl_black_box_vo_net;
  o_re_2 <= reinterpret25_output_port_net;
  o_re_3 <= reinterpret26_output_port_net;
  o_re_4 <= reinterpret27_output_port_net;
  o_re_5 <= reinterpret28_output_port_net;
  o_re_6 <= reinterpret29_output_port_net;
  o_re_7 <= reinterpret30_output_port_net;
  o_re_8 <= reinterpret31_output_port_net;
  o_im_2 <= reinterpret17_output_port_net;
  o_im_3 <= reinterpret18_output_port_net;
  o_im_4 <= reinterpret19_output_port_net;
  o_im_5 <= reinterpret20_output_port_net;
  o_im_6 <= reinterpret21_output_port_net;
  o_im_7 <= reinterpret22_output_port_net;
  o_im_8 <= reinterpret23_output_port_net;
  mux2_y_net <= i_re_1;
  mux27_y_net <= i_im_1;
  delay11_q_net <= vi;
  constant15_op_net <= si;
  mux29_y_net <= i_re_2;
  mux33_y_net <= i_re_3;
  mux37_y_net <= i_re_4;
  mux41_y_net <= i_re_5;
  mux45_y_net <= i_re_6;
  mux49_y_net <= i_re_7;
  mux53_y_net <= i_re_8;
  mux30_y_net <= i_im_2;
  mux34_y_net <= i_im_3;
  mux38_y_net <= i_im_4;
  mux42_y_net <= i_im_5;
  mux46_y_net <= i_im_6;
  mux50_y_net <= i_im_7;
  mux54_y_net <= i_im_8;
  clk_net <= clk_1;
  ce_net <= ce_1;
  vector_fft : entity xil_defaultlib.psb3_0_vector_fft 
  port map (
    i_re_1 => mux27_y_net,
    i_im_1 => mux2_y_net,
    vi => delay11_q_net,
    si => constant15_op_net,
    i_re_2 => mux30_y_net,
    i_re_3 => mux34_y_net,
    i_re_4 => mux38_y_net,
    i_re_5 => mux42_y_net,
    i_re_6 => mux46_y_net,
    i_re_7 => mux50_y_net,
    i_re_8 => mux54_y_net,
    i_im_2 => mux29_y_net,
    i_im_3 => mux33_y_net,
    i_im_4 => mux37_y_net,
    i_im_5 => mux41_y_net,
    i_im_6 => mux45_y_net,
    i_im_7 => mux49_y_net,
    i_im_8 => mux53_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    o_re_1 => reinterpret16_output_port_net,
    o_im_1 => reinterpret24_output_port_net,
    vo => test_systolicfft_vhdl_black_box_vo_net,
    o_re_2 => reinterpret17_output_port_net,
    o_re_3 => reinterpret18_output_port_net,
    o_re_4 => reinterpret19_output_port_net,
    o_re_5 => reinterpret20_output_port_net,
    o_re_6 => reinterpret21_output_port_net,
    o_re_7 => reinterpret22_output_port_net,
    o_re_8 => reinterpret23_output_port_net,
    o_im_2 => reinterpret25_output_port_net,
    o_im_3 => reinterpret26_output_port_net,
    o_im_4 => reinterpret27_output_port_net,
    o_im_5 => reinterpret28_output_port_net,
    o_im_6 => reinterpret29_output_port_net,
    o_im_7 => reinterpret30_output_port_net,
    o_im_8 => reinterpret31_output_port_net
  );
end structural;
-- Generated from Simulink block PSB3_0_struct
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_struct is
  port (
    gin_tl_reset : in std_logic_vector( 1-1 downto 0 );
    gin_tl_start : in std_logic_vector( 1-1 downto 0 );
    gin_addr : in std_logic_vector( 8-1 downto 0 );
    gin_dphi : in std_logic_vector( 16-1 downto 0 );
    gin_init_im : in std_logic_vector( 18-1 downto 0 );
    gin_init_re : in std_logic_vector( 18-1 downto 0 );
    gin_we_even_1 : in std_logic_vector( 1-1 downto 0 );
    gin_we_even_2 : in std_logic_vector( 1-1 downto 0 );
    gin_we_even_3 : in std_logic_vector( 1-1 downto 0 );
    gin_we_even_4 : in std_logic_vector( 1-1 downto 0 );
    gin_we_odd_1 : in std_logic_vector( 1-1 downto 0 );
    gin_we_odd_2 : in std_logic_vector( 1-1 downto 0 );
    gin_we_odd_3 : in std_logic_vector( 1-1 downto 0 );
    gin_we_odd_4 : in std_logic_vector( 1-1 downto 0 );
    ts_0 : in std_logic_vector( 12-1 downto 0 );
    ts_1 : in std_logic_vector( 12-1 downto 0 );
    ts_2 : in std_logic_vector( 12-1 downto 0 );
    ts_3 : in std_logic_vector( 12-1 downto 0 );
    ts_4 : in std_logic_vector( 12-1 downto 0 );
    ts_5 : in std_logic_vector( 12-1 downto 0 );
    ts_6 : in std_logic_vector( 12-1 downto 0 );
    ts_7 : in std_logic_vector( 12-1 downto 0 );
    ts_a : in std_logic_vector( 8-1 downto 0 );
    ts_w : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    gout_cordic_delay_even_1 : out std_logic_vector( 12-1 downto 0 );
    gout_psb_tvalid : out std_logic_vector( 1-1 downto 0 );
    gout_delay_ifft : out std_logic_vector( 12-1 downto 0 );
    gout_ov_ifft : out std_logic_vector( 1-1 downto 0 );
    gout_ov_add : out std_logic_vector( 1-1 downto 0 );
    gout_psb_im_0 : out std_logic_vector( 16-1 downto 0 );
    gout_psb_im_1 : out std_logic_vector( 16-1 downto 0 );
    gout_psb_im_2 : out std_logic_vector( 16-1 downto 0 );
    gout_psb_im_3 : out std_logic_vector( 16-1 downto 0 );
    gout_psb_re_0 : out std_logic_vector( 16-1 downto 0 );
    gout_psb_re_1 : out std_logic_vector( 16-1 downto 0 );
    gout_psb_re_2 : out std_logic_vector( 16-1 downto 0 );
    gout_psb_re_3 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0_struct;
architecture structural of psb3_0_struct is 
  signal gin_addr_net : std_logic_vector( 8-1 downto 0 );
  signal gin_tl_reset_net : std_logic_vector( 1-1 downto 0 );
  signal gin_tl_start_net : std_logic_vector( 1-1 downto 0 );
  signal expression1_dout_net : std_logic_vector( 1-1 downto 0 );
  signal ts_1_net : std_logic_vector( 12-1 downto 0 );
  signal ts_2_net : std_logic_vector( 12-1 downto 0 );
  signal gin_we_odd_2_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret6_output_port_net_x14 : std_logic_vector( 16-1 downto 0 );
  signal gin_we_even_2_net : std_logic_vector( 1-1 downto 0 );
  signal expression_dout_net : std_logic_vector( 1-1 downto 0 );
  signal ts_a_net : std_logic_vector( 8-1 downto 0 );
  signal gin_we_odd_4_net : std_logic_vector( 1-1 downto 0 );
  signal ts_w_net : std_logic_vector( 1-1 downto 0 );
  signal counter1_op_net_x7 : std_logic_vector( 12-1 downto 0 );
  signal ts_6_net : std_logic_vector( 12-1 downto 0 );
  signal reinterpret2_output_port_net_x14 : std_logic_vector( 16-1 downto 0 );
  signal ts_5_net : std_logic_vector( 12-1 downto 0 );
  signal reinterpret1_output_port_net_x14 : std_logic_vector( 16-1 downto 0 );
  signal ts_0_net : std_logic_vector( 12-1 downto 0 );
  signal gin_init_im_net : std_logic_vector( 18-1 downto 0 );
  signal ts_7_net : std_logic_vector( 12-1 downto 0 );
  signal gin_we_even_4_net : std_logic_vector( 1-1 downto 0 );
  signal counter1_op_net_x6 : std_logic_vector( 12-1 downto 0 );
  signal ts_3_net : std_logic_vector( 12-1 downto 0 );
  signal ts_4_net : std_logic_vector( 12-1 downto 0 );
  signal reinterpret3_output_port_net_x14 : std_logic_vector( 16-1 downto 0 );
  signal gin_we_odd_3_net : std_logic_vector( 1-1 downto 0 );
  signal gin_we_odd_1_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret7_output_port_net_x14 : std_logic_vector( 16-1 downto 0 );
  signal gin_dphi_net : std_logic_vector( 16-1 downto 0 );
  signal gin_init_re_net : std_logic_vector( 18-1 downto 0 );
  signal gin_we_even_1_net : std_logic_vector( 1-1 downto 0 );
  signal gin_we_even_3_net : std_logic_vector( 1-1 downto 0 );
  signal delay54_q_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net_x17 : std_logic_vector( 16-1 downto 0 );
  signal clk_net : std_logic;
  signal delay37_q_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net_x18 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net_x17 : std_logic_vector( 16-1 downto 0 );
  signal delay48_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret0_output_port_net_x16 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net_x17 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net_x14 : std_logic_vector( 16-1 downto 0 );
  signal cordic_6_0_even_1_m_axis_dout_tdata_imag_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal cordic_6_0_even_2_m_axis_dout_tdata_real_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net_x18 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net_x18 : std_logic_vector( 16-1 downto 0 );
  signal delay31_q_net : std_logic_vector( 1-1 downto 0 );
  signal cordic_6_0_even_2_m_axis_dout_tdata_real_net : std_logic_vector( 16-1 downto 0 );
  signal cordic_6_0_odd_2_m_axis_dout_tdata_real_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net_x18 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net_x18 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net_x17 : std_logic_vector( 16-1 downto 0 );
  signal delay44_q_net : std_logic_vector( 18-1 downto 0 );
  signal cordic_6_0_odd_1_m_axis_dout_tdata_real_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net_x17 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net_x17 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net_x17 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net_x14 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net_x17 : std_logic_vector( 16-1 downto 0 );
  signal delay8_q_net_x3 : std_logic_vector( 1-1 downto 0 );
  signal delay38_q_net : std_logic_vector( 8-1 downto 0 );
  signal register_q_net_x7 : std_logic_vector( 1-1 downto 0 );
  signal reinterpret4_output_port_net_x17 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net_x17 : std_logic_vector( 16-1 downto 0 );
  signal cordic_6_0_odd_1_m_axis_dout_tdata_imag_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal cordic_6_0_even_1_m_axis_dout_tdata_real_net : std_logic_vector( 16-1 downto 0 );
  signal cordic_6_0_even_2_m_axis_dout_tdata_imag_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net_x18 : std_logic_vector( 16-1 downto 0 );
  signal ram_dphi_addr_op_net : std_logic_vector( 8-1 downto 0 );
  signal cordic_6_0_even_1_m_axis_dout_tdata_imag_net : std_logic_vector( 16-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal cordic_6_0_odd_1_m_axis_dout_tdata_imag_net : std_logic_vector( 16-1 downto 0 );
  signal ce_net : std_logic;
  signal cordic_6_0_odd_2_m_axis_dout_tdata_imag_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net_x18 : std_logic_vector( 16-1 downto 0 );
  signal delay35_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay49_q_net : std_logic_vector( 1-1 downto 0 );
  signal cordic_6_0_odd_2_m_axis_dout_tdata_real_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal delay43_q_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret1_output_port_net_x17 : std_logic_vector( 16-1 downto 0 );
  signal delay14_q_net : std_logic_vector( 1-1 downto 0 );
  signal cordic_6_0_odd_1_m_axis_dout_tdata_real_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net_x17 : std_logic_vector( 16-1 downto 0 );
  signal cordic_6_0_even_1_m_axis_dout_tdata_real_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal cordic_6_0_even_2_m_axis_dout_tdata_imag_net : std_logic_vector( 16-1 downto 0 );
  signal cordic_6_0_even_1_m_axis_dout_tvalid_net_x0 : std_logic;
  signal cordic_6_0_odd_2_m_axis_dout_tdata_imag_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net_x17 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net_x17 : std_logic_vector( 16-1 downto 0 );
  signal delay26_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret0_output_port_net_x17 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net_x18 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net_x15 : std_logic_vector( 16-1 downto 0 );
  signal addsub0_s_net_x5 : std_logic_vector( 16-1 downto 0 );
  signal mult0_p_net_x6 : std_logic_vector( 16-1 downto 0 );
  signal mult4_p_net_x6 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net_x16 : std_logic_vector( 16-1 downto 0 );
  signal mult7_p_net_x6 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net_x15 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net_x16 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net_x14 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net_x16 : std_logic_vector( 16-1 downto 0 );
  signal mult8_p_net_x6 : std_logic_vector( 16-1 downto 0 );
  signal mult9_p_net_x6 : std_logic_vector( 16-1 downto 0 );
  signal mult12_p_net_x6 : std_logic_vector( 16-1 downto 0 );
  signal mult13_p_net_x6 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net_x15 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net_x16 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net_x15 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net_x15 : std_logic_vector( 16-1 downto 0 );
  signal mult14_p_net_x6 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net_x14 : std_logic_vector( 16-1 downto 0 );
  signal mult15_p_net_x6 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net_x16 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net_x4 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net_x16 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net_x15 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net_x15 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net_x14 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net_x16 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net_x15 : std_logic_vector( 16-1 downto 0 );
  signal register_q_net_x6 : std_logic_vector( 1-1 downto 0 );
  signal mult1_p_net_x6 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net_x17 : std_logic_vector( 16-1 downto 0 );
  signal mult3_p_net_x6 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net_x15 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net_x15 : std_logic_vector( 16-1 downto 0 );
  signal mult6_p_net_x6 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net_x16 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net_x14 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net_x15 : std_logic_vector( 16-1 downto 0 );
  signal mult10_p_net_x6 : std_logic_vector( 16-1 downto 0 );
  signal mult11_p_net_x6 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net_x4 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net_x4 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net_x14 : std_logic_vector( 16-1 downto 0 );
  signal mult5_p_net_x6 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net_x16 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net_x16 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net_x16 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net_x15 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net_x14 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net_x15 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net_x14 : std_logic_vector( 16-1 downto 0 );
  signal mult2_p_net_x6 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net_x16 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net_x16 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net_x16 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net_x15 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net_x16 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net_x15 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net_x15 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net_x14 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net_x4 : std_logic_vector( 16-1 downto 0 );
  signal fifo6_full_net : std_logic;
  signal fifo3_full_net : std_logic;
  signal fifo5_empty_net : std_logic;
  signal fifo4_empty_net : std_logic;
  signal fifo2_full_net : std_logic;
  signal fifo4_full_net : std_logic;
  signal fifo3_empty_net : std_logic;
  signal fifo6_empty_net : std_logic;
  signal fifo2_empty_net : std_logic;
  signal fifo5_full_net : std_logic;
  signal reinterpret3_output_port_net_x1 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net_x1 : std_logic_vector( 16-1 downto 0 );
  signal addsub10_s_net_x5 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net_x4 : std_logic_vector( 16-1 downto 0 );
  signal addsub2_s_net_x5 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net_x1 : std_logic_vector( 16-1 downto 0 );
  signal addsub4_s_net_x5 : std_logic_vector( 16-1 downto 0 );
  signal addsub5_s_net_x5 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net_x1 : std_logic_vector( 16-1 downto 0 );
  signal mult12_p_net_x5 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net_x1 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net_x4 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net_x4 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net_x1 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net_x1 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net_x1 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net_x4 : std_logic_vector( 16-1 downto 0 );
  signal addsub15_s_net_x5 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net_x1 : std_logic_vector( 16-1 downto 0 );
  signal mult2_p_net_x5 : std_logic_vector( 16-1 downto 0 );
  signal addsub7_s_net_x5 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net_x1 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net_x1 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net_x1 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net_x1 : std_logic_vector( 16-1 downto 0 );
  signal addsub0_s_net_x3 : std_logic_vector( 16-1 downto 0 );
  signal mult8_p_net_x5 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net_x4 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net_x1 : std_logic_vector( 16-1 downto 0 );
  signal mult10_p_net_x5 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net_x4 : std_logic_vector( 16-1 downto 0 );
  signal addsub6_s_net_x4 : std_logic_vector( 16-1 downto 0 );
  signal addsub1_s_net_x3 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net_x4 : std_logic_vector( 16-1 downto 0 );
  signal addsub2_s_net_x3 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net_x1 : std_logic_vector( 16-1 downto 0 );
  signal addsub3_s_net_x3 : std_logic_vector( 16-1 downto 0 );
  signal addsub13_s_net_x5 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net_x1 : std_logic_vector( 16-1 downto 0 );
  signal mult9_p_net_x5 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net_x4 : std_logic_vector( 16-1 downto 0 );
  signal addsub8_s_net_x5 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net_x4 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net_x4 : std_logic_vector( 16-1 downto 0 );
  signal register_q_net_x5 : std_logic_vector( 1-1 downto 0 );
  signal addsub11_s_net_x5 : std_logic_vector( 16-1 downto 0 );
  signal addsub9_s_net_x5 : std_logic_vector( 16-1 downto 0 );
  signal mult1_p_net_x5 : std_logic_vector( 16-1 downto 0 );
  signal addsub14_s_net_x5 : std_logic_vector( 16-1 downto 0 );
  signal mult3_p_net_x5 : std_logic_vector( 16-1 downto 0 );
  signal mult4_p_net_x5 : std_logic_vector( 16-1 downto 0 );
  signal mult5_p_net_x5 : std_logic_vector( 16-1 downto 0 );
  signal mult0_p_net_x5 : std_logic_vector( 16-1 downto 0 );
  signal addsub3_s_net_x5 : std_logic_vector( 16-1 downto 0 );
  signal mult6_p_net_x5 : std_logic_vector( 16-1 downto 0 );
  signal mult7_p_net_x5 : std_logic_vector( 16-1 downto 0 );
  signal mult11_p_net_x5 : std_logic_vector( 16-1 downto 0 );
  signal addsub12_s_net_x5 : std_logic_vector( 16-1 downto 0 );
  signal mult13_p_net_x5 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net_x4 : std_logic_vector( 16-1 downto 0 );
  signal mult14_p_net_x5 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net_x4 : std_logic_vector( 16-1 downto 0 );
  signal addsub1_s_net_x5 : std_logic_vector( 16-1 downto 0 );
  signal mult15_p_net_x5 : std_logic_vector( 16-1 downto 0 );
  signal addsub6_s_net_x2 : std_logic_vector( 16-1 downto 0 );
  signal mult11_p_net_x4 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net_x11 : std_logic_vector( 16-1 downto 0 );
  signal addsub14_s_net_x1 : std_logic_vector( 16-1 downto 0 );
  signal mult5_p_net_x4 : std_logic_vector( 16-1 downto 0 );
  signal mult9_p_net_x4 : std_logic_vector( 16-1 downto 0 );
  signal addsub10_s_net_x1 : std_logic_vector( 16-1 downto 0 );
  signal addsub2_s_net_x1 : std_logic_vector( 16-1 downto 0 );
  signal addsub0_s_net_x1 : std_logic_vector( 16-1 downto 0 );
  signal addsub9_s_net_x3 : std_logic_vector( 16-1 downto 0 );
  signal addsub8_s_net_x3 : std_logic_vector( 16-1 downto 0 );
  signal mult10_p_net_x4 : std_logic_vector( 16-1 downto 0 );
  signal addsub10_s_net_x3 : std_logic_vector( 16-1 downto 0 );
  signal addsub5_s_net_x3 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net_x11 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net_x11 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net_x11 : std_logic_vector( 16-1 downto 0 );
  signal mult8_p_net_x4 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net_x11 : std_logic_vector( 16-1 downto 0 );
  signal addsub11_s_net_x1 : std_logic_vector( 16-1 downto 0 );
  signal mult0_p_net_x4 : std_logic_vector( 16-1 downto 0 );
  signal addsub13_s_net_x1 : std_logic_vector( 16-1 downto 0 );
  signal mult13_p_net_x4 : std_logic_vector( 16-1 downto 0 );
  signal addsub15_s_net_x1 : std_logic_vector( 16-1 downto 0 );
  signal mult14_p_net_x4 : std_logic_vector( 16-1 downto 0 );
  signal register_q_net_x3 : std_logic_vector( 1-1 downto 0 );
  signal addsub4_s_net_x3 : std_logic_vector( 16-1 downto 0 );
  signal addsub12_s_net_x3 : std_logic_vector( 16-1 downto 0 );
  signal mult1_p_net_x4 : std_logic_vector( 16-1 downto 0 );
  signal addsub7_s_net_x1 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net_x11 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net_x11 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net_x11 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net_x11 : std_logic_vector( 16-1 downto 0 );
  signal addsub1_s_net_x1 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net_x11 : std_logic_vector( 16-1 downto 0 );
  signal addsub12_s_net_x1 : std_logic_vector( 16-1 downto 0 );
  signal mult0_p_net_x3 : std_logic_vector( 16-1 downto 0 );
  signal mult12_p_net_x4 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net_x8 : std_logic_vector( 16-1 downto 0 );
  signal register_q_net_x4 : std_logic_vector( 1-1 downto 0 );
  signal addsub15_s_net_x3 : std_logic_vector( 16-1 downto 0 );
  signal mult15_p_net_x4 : std_logic_vector( 16-1 downto 0 );
  signal addsub13_s_net_x3 : std_logic_vector( 16-1 downto 0 );
  signal addsub14_s_net_x3 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net_x11 : std_logic_vector( 16-1 downto 0 );
  signal addsub11_s_net_x3 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net_x11 : std_logic_vector( 16-1 downto 0 );
  signal mult2_p_net_x4 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net_x11 : std_logic_vector( 16-1 downto 0 );
  signal mult3_p_net_x4 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net_x11 : std_logic_vector( 16-1 downto 0 );
  signal addsub4_s_net_x1 : std_logic_vector( 16-1 downto 0 );
  signal mult6_p_net_x4 : std_logic_vector( 16-1 downto 0 );
  signal addsub3_s_net_x1 : std_logic_vector( 16-1 downto 0 );
  signal mult7_p_net_x4 : std_logic_vector( 16-1 downto 0 );
  signal addsub5_s_net_x1 : std_logic_vector( 16-1 downto 0 );
  signal addsub6_s_net_x6 : std_logic_vector( 16-1 downto 0 );
  signal addsub8_s_net_x1 : std_logic_vector( 16-1 downto 0 );
  signal addsub9_s_net_x1 : std_logic_vector( 16-1 downto 0 );
  signal addsub7_s_net_x3 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net_x11 : std_logic_vector( 16-1 downto 0 );
  signal mult4_p_net_x4 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net_x11 : std_logic_vector( 16-1 downto 0 );
  signal mult6_p_net_x3 : std_logic_vector( 16-1 downto 0 );
  signal addsub14_s_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net_x8 : std_logic_vector( 16-1 downto 0 );
  signal addsub15_s_net : std_logic_vector( 16-1 downto 0 );
  signal mult0_p_net_x2 : std_logic_vector( 16-1 downto 0 );
  signal mult2_p_net_x2 : std_logic_vector( 16-1 downto 0 );
  signal addsub8_s_net : std_logic_vector( 16-1 downto 0 );
  signal mult4_p_net_x2 : std_logic_vector( 16-1 downto 0 );
  signal mult7_p_net_x2 : std_logic_vector( 16-1 downto 0 );
  signal mult7_p_net_x3 : std_logic_vector( 16-1 downto 0 );
  signal register_q_net_x2 : std_logic_vector( 1-1 downto 0 );
  signal mult5_p_net_x2 : std_logic_vector( 16-1 downto 0 );
  signal mult6_p_net_x2 : std_logic_vector( 16-1 downto 0 );
  signal mult8_p_net_x2 : std_logic_vector( 16-1 downto 0 );
  signal mult9_p_net_x2 : std_logic_vector( 16-1 downto 0 );
  signal addsub0_s_net_x6 : std_logic_vector( 16-1 downto 0 );
  signal mult10_p_net_x2 : std_logic_vector( 16-1 downto 0 );
  signal mult12_p_net_x2 : std_logic_vector( 16-1 downto 0 );
  signal mult14_p_net_x2 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net_x8 : std_logic_vector( 16-1 downto 0 );
  signal mult12_p_net_x3 : std_logic_vector( 16-1 downto 0 );
  signal mult3_p_net_x2 : std_logic_vector( 16-1 downto 0 );
  signal mult13_p_net_x2 : std_logic_vector( 16-1 downto 0 );
  signal mult2_p_net_x3 : std_logic_vector( 16-1 downto 0 );
  signal addsub0_s_net : std_logic_vector( 16-1 downto 0 );
  signal mult11_p_net_x3 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net_x8 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net_x5 : std_logic_vector( 16-1 downto 0 );
  signal addsub13_s_net : std_logic_vector( 16-1 downto 0 );
  signal mult5_p_net_x3 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net_x8 : std_logic_vector( 16-1 downto 0 );
  signal mult1_p_net_x2 : std_logic_vector( 16-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 16-1 downto 0 );
  signal mult11_p_net_x2 : std_logic_vector( 16-1 downto 0 );
  signal addsub5_s_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net_x8 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net_x8 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net_x8 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net_x8 : std_logic_vector( 16-1 downto 0 );
  signal mult4_p_net_x3 : std_logic_vector( 16-1 downto 0 );
  signal mult10_p_net_x3 : std_logic_vector( 16-1 downto 0 );
  signal mult8_p_net_x3 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net_x8 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net_x8 : std_logic_vector( 16-1 downto 0 );
  signal mult1_p_net_x3 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net_x8 : std_logic_vector( 16-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub9_s_net : std_logic_vector( 16-1 downto 0 );
  signal mult13_p_net_x3 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net_x8 : std_logic_vector( 16-1 downto 0 );
  signal mult15_p_net_x3 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net_x8 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net_x8 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net_x8 : std_logic_vector( 16-1 downto 0 );
  signal mult9_p_net_x3 : std_logic_vector( 16-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub10_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub11_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub12_s_net : std_logic_vector( 16-1 downto 0 );
  signal mult3_p_net_x3 : std_logic_vector( 16-1 downto 0 );
  signal mult14_p_net_x3 : std_logic_vector( 16-1 downto 0 );
  signal addsub3_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub6_s_net : std_logic_vector( 16-1 downto 0 );
  signal addsub7_s_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net_x5 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net_x5 : std_logic_vector( 16-1 downto 0 );
  signal mult2_p_net_x1 : std_logic_vector( 16-1 downto 0 );
  signal mult8_p_net_x1 : std_logic_vector( 16-1 downto 0 );
  signal mult1_p_net_x1 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net_x13 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net_x5 : std_logic_vector( 16-1 downto 0 );
  signal mult13_p_net_x1 : std_logic_vector( 16-1 downto 0 );
  signal mult4_p_net_x1 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net_x5 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net_x5 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net_x13 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net_x5 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net_x5 : std_logic_vector( 16-1 downto 0 );
  signal addsub1_s_net_x6 : std_logic_vector( 16-1 downto 0 );
  signal addsub14_s_net_x6 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net_x13 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net_x13 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net_x13 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net_x5 : std_logic_vector( 16-1 downto 0 );
  signal addsub11_s_net_x6 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net_x13 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net_x5 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net_x13 : std_logic_vector( 16-1 downto 0 );
  signal register_q_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal reinterpret4_output_port_net_x5 : std_logic_vector( 16-1 downto 0 );
  signal addsub3_s_net_x6 : std_logic_vector( 16-1 downto 0 );
  signal addsub12_s_net_x6 : std_logic_vector( 16-1 downto 0 );
  signal addsub10_s_net_x6 : std_logic_vector( 16-1 downto 0 );
  signal addsub0_s_net_x4 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net_x13 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net_x13 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net_x13 : std_logic_vector( 16-1 downto 0 );
  signal mult12_p_net_x1 : std_logic_vector( 16-1 downto 0 );
  signal mult10_p_net_x1 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net_x13 : std_logic_vector( 16-1 downto 0 );
  signal addsub9_s_net_x6 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net_x13 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net_x13 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net_x5 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net_x13 : std_logic_vector( 16-1 downto 0 );
  signal addsub6_s_net_x5 : std_logic_vector( 16-1 downto 0 );
  signal addsub15_s_net_x6 : std_logic_vector( 16-1 downto 0 );
  signal addsub4_s_net_x6 : std_logic_vector( 16-1 downto 0 );
  signal addsub5_s_net_x6 : std_logic_vector( 16-1 downto 0 );
  signal mult7_p_net_x1 : std_logic_vector( 16-1 downto 0 );
  signal addsub2_s_net_x6 : std_logic_vector( 16-1 downto 0 );
  signal mult11_p_net_x1 : std_logic_vector( 16-1 downto 0 );
  signal mult15_p_net_x1 : std_logic_vector( 16-1 downto 0 );
  signal mult0_p_net_x1 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net_x13 : std_logic_vector( 16-1 downto 0 );
  signal mult6_p_net_x1 : std_logic_vector( 16-1 downto 0 );
  signal mult15_p_net_x2 : std_logic_vector( 16-1 downto 0 );
  signal addsub13_s_net_x6 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net_x5 : std_logic_vector( 16-1 downto 0 );
  signal mult9_p_net_x1 : std_logic_vector( 16-1 downto 0 );
  signal mult5_p_net_x1 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net_x5 : std_logic_vector( 16-1 downto 0 );
  signal mult14_p_net_x1 : std_logic_vector( 16-1 downto 0 );
  signal addsub8_s_net_x6 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net_x5 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net_x5 : std_logic_vector( 16-1 downto 0 );
  signal addsub7_s_net_x6 : std_logic_vector( 16-1 downto 0 );
  signal mult3_p_net_x1 : std_logic_vector( 16-1 downto 0 );
  signal mult11_p_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net_x12 : std_logic_vector( 16-1 downto 0 );
  signal addsub6_s_net_x3 : std_logic_vector( 16-1 downto 0 );
  signal addsub10_s_net_x4 : std_logic_vector( 16-1 downto 0 );
  signal mult3_p_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net_x12 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net_x12 : std_logic_vector( 16-1 downto 0 );
  signal mult14_p_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net_x12 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net_x12 : std_logic_vector( 16-1 downto 0 );
  signal mult0_p_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal register_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal reinterpret13_output_port_net_x12 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net_x12 : std_logic_vector( 16-1 downto 0 );
  signal addsub2_s_net_x2 : std_logic_vector( 16-1 downto 0 );
  signal addsub5_s_net_x2 : std_logic_vector( 16-1 downto 0 );
  signal addsub2_s_net_x4 : std_logic_vector( 16-1 downto 0 );
  signal mult6_p_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net_x12 : std_logic_vector( 16-1 downto 0 );
  signal addsub3_s_net_x2 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net_x12 : std_logic_vector( 16-1 downto 0 );
  signal addsub7_s_net_x2 : std_logic_vector( 16-1 downto 0 );
  signal addsub9_s_net_x2 : std_logic_vector( 16-1 downto 0 );
  signal addsub8_s_net_x2 : std_logic_vector( 16-1 downto 0 );
  signal addsub12_s_net_x2 : std_logic_vector( 16-1 downto 0 );
  signal addsub5_s_net_x4 : std_logic_vector( 16-1 downto 0 );
  signal addsub12_s_net_x4 : std_logic_vector( 16-1 downto 0 );
  signal addsub3_s_net_x4 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net_x12 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net_x12 : std_logic_vector( 16-1 downto 0 );
  signal addsub4_s_net_x2 : std_logic_vector( 16-1 downto 0 );
  signal addsub6_s_net_x1 : std_logic_vector( 16-1 downto 0 );
  signal addsub13_s_net_x4 : std_logic_vector( 16-1 downto 0 );
  signal mult13_p_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal addsub11_s_net_x2 : std_logic_vector( 16-1 downto 0 );
  signal addsub13_s_net_x2 : std_logic_vector( 16-1 downto 0 );
  signal addsub14_s_net_x2 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net_x13 : std_logic_vector( 16-1 downto 0 );
  signal addsub9_s_net_x4 : std_logic_vector( 16-1 downto 0 );
  signal addsub1_s_net_x2 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net_x12 : std_logic_vector( 16-1 downto 0 );
  signal addsub10_s_net_x2 : std_logic_vector( 16-1 downto 0 );
  signal addsub11_s_net_x4 : std_logic_vector( 16-1 downto 0 );
  signal addsub14_s_net_x4 : std_logic_vector( 16-1 downto 0 );
  signal mult12_p_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal addsub7_s_net_x4 : std_logic_vector( 16-1 downto 0 );
  signal mult4_p_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal addsub0_s_net_x2 : std_logic_vector( 16-1 downto 0 );
  signal addsub1_s_net_x4 : std_logic_vector( 16-1 downto 0 );
  signal mult8_p_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal mult1_p_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net_x12 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net_x12 : std_logic_vector( 16-1 downto 0 );
  signal mult7_p_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal addsub4_s_net_x4 : std_logic_vector( 16-1 downto 0 );
  signal mult5_p_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net_x12 : std_logic_vector( 16-1 downto 0 );
  signal addsub8_s_net_x4 : std_logic_vector( 16-1 downto 0 );
  signal mult10_p_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal mult15_p_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net_x12 : std_logic_vector( 16-1 downto 0 );
  signal addsub15_s_net_x4 : std_logic_vector( 16-1 downto 0 );
  signal mult2_p_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal mult9_p_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal slice1_y_net_x6 : std_logic_vector( 16-1 downto 0 );
  signal slice2_y_net_x6 : std_logic_vector( 16-1 downto 0 );
  signal slice3_y_net_x6 : std_logic_vector( 16-1 downto 0 );
  signal slice4_y_net_x6 : std_logic_vector( 16-1 downto 0 );
  signal slice5_y_net_x6 : std_logic_vector( 16-1 downto 0 );
  signal slice6_y_net_x6 : std_logic_vector( 16-1 downto 0 );
  signal addsub12_s_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal slice7_y_net_x6 : std_logic_vector( 16-1 downto 0 );
  signal mult1_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net_x26 : std_logic_vector( 16-1 downto 0 );
  signal addsub8_s_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal slice8_y_net_x6 : std_logic_vector( 16-1 downto 0 );
  signal mult3_p_net : std_logic_vector( 16-1 downto 0 );
  signal slice9_y_net_x6 : std_logic_vector( 16-1 downto 0 );
  signal addsub15_s_net_x2 : std_logic_vector( 16-1 downto 0 );
  signal addsub13_s_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal slice10_y_net_x6 : std_logic_vector( 16-1 downto 0 );
  signal slice11_y_net_x6 : std_logic_vector( 16-1 downto 0 );
  signal slice12_y_net_x6 : std_logic_vector( 16-1 downto 0 );
  signal mult5_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult14_p_net : std_logic_vector( 16-1 downto 0 );
  signal slice13_y_net_x6 : std_logic_vector( 16-1 downto 0 );
  signal addsub0_s_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal addsub1_s_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal addsub10_s_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net_x26 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net_x26 : std_logic_vector( 16-1 downto 0 );
  signal mult11_p_net : std_logic_vector( 16-1 downto 0 );
  signal addsub9_s_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net_x27 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net_x26 : std_logic_vector( 16-1 downto 0 );
  signal addsub4_s_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal addsub5_s_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal addsub7_s_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal addsub11_s_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal mult12_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult6_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult15_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult9_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net_x27 : std_logic_vector( 16-1 downto 0 );
  signal mult0_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult2_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult10_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net_x27 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net_x27 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net_x26 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net_x26 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net_x26 : std_logic_vector( 16-1 downto 0 );
  signal register_q_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret7_output_port_net_x27 : std_logic_vector( 16-1 downto 0 );
  signal addsub2_s_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal addsub3_s_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal mult4_p_net : std_logic_vector( 16-1 downto 0 );
  signal mult13_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net_x26 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net_x26 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net_x27 : std_logic_vector( 16-1 downto 0 );
  signal addsub6_s_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal mult7_p_net : std_logic_vector( 16-1 downto 0 );
  signal addsub14_s_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal addsub15_s_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal mult8_p_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net_x27 : std_logic_vector( 16-1 downto 0 );
  signal slice0_y_net_x6 : std_logic_vector( 16-1 downto 0 );
  signal slice2_y_net_x4 : std_logic_vector( 16-1 downto 0 );
  signal slice12_y_net_x3 : std_logic_vector( 16-1 downto 0 );
  signal slice6_y_net_x2 : std_logic_vector( 16-1 downto 0 );
  signal slice7_y_net_x2 : std_logic_vector( 16-1 downto 0 );
  signal slice9_y_net_x4 : std_logic_vector( 16-1 downto 0 );
  signal slice13_y_net_x4 : std_logic_vector( 16-1 downto 0 );
  signal bitbasher1_a_net : std_logic_vector( 256-1 downto 0 );
  signal slice8_y_net_x4 : std_logic_vector( 16-1 downto 0 );
  signal slice1_y_net_x3 : std_logic_vector( 16-1 downto 0 );
  signal slice7_y_net_x3 : std_logic_vector( 16-1 downto 0 );
  signal slice8_y_net_x3 : std_logic_vector( 16-1 downto 0 );
  signal slice6_y_net_x5 : std_logic_vector( 16-1 downto 0 );
  signal slice4_y_net_x5 : std_logic_vector( 16-1 downto 0 );
  signal slice15_y_net_x5 : std_logic_vector( 16-1 downto 0 );
  signal slice3_y_net_x4 : std_logic_vector( 16-1 downto 0 );
  signal slice9_y_net_x5 : std_logic_vector( 16-1 downto 0 );
  signal slice5_y_net_x4 : std_logic_vector( 16-1 downto 0 );
  signal slice6_y_net_x3 : std_logic_vector( 16-1 downto 0 );
  signal slice1_y_net_x2 : std_logic_vector( 16-1 downto 0 );
  signal slice8_y_net_x5 : std_logic_vector( 16-1 downto 0 );
  signal bitbasher2_a_net : std_logic_vector( 256-1 downto 0 );
  signal slice15_y_net_x4 : std_logic_vector( 16-1 downto 0 );
  signal slice2_y_net_x2 : std_logic_vector( 16-1 downto 0 );
  signal slice8_y_net_x2 : std_logic_vector( 16-1 downto 0 );
  signal slice9_y_net_x2 : std_logic_vector( 16-1 downto 0 );
  signal slice10_y_net_x5 : std_logic_vector( 16-1 downto 0 );
  signal slice2_y_net_x5 : std_logic_vector( 16-1 downto 0 );
  signal slice9_y_net_x3 : std_logic_vector( 16-1 downto 0 );
  signal slice11_y_net_x4 : std_logic_vector( 16-1 downto 0 );
  signal slice1_y_net_x4 : std_logic_vector( 16-1 downto 0 );
  signal slice11_y_net_x5 : std_logic_vector( 16-1 downto 0 );
  signal slice11_y_net_x3 : std_logic_vector( 16-1 downto 0 );
  signal slice2_y_net_x3 : std_logic_vector( 16-1 downto 0 );
  signal slice10_y_net_x3 : std_logic_vector( 16-1 downto 0 );
  signal slice15_y_net_x3 : std_logic_vector( 16-1 downto 0 );
  signal slice0_y_net_x2 : std_logic_vector( 16-1 downto 0 );
  signal slice3_y_net_x3 : std_logic_vector( 16-1 downto 0 );
  signal slice4_y_net_x4 : std_logic_vector( 16-1 downto 0 );
  signal slice4_y_net_x3 : std_logic_vector( 16-1 downto 0 );
  signal slice0_y_net_x4 : std_logic_vector( 16-1 downto 0 );
  signal slice3_y_net_x2 : std_logic_vector( 16-1 downto 0 );
  signal slice5_y_net_x5 : std_logic_vector( 16-1 downto 0 );
  signal slice7_y_net_x5 : std_logic_vector( 16-1 downto 0 );
  signal slice14_y_net_x6 : std_logic_vector( 16-1 downto 0 );
  signal slice13_y_net_x5 : std_logic_vector( 16-1 downto 0 );
  signal slice6_y_net_x4 : std_logic_vector( 16-1 downto 0 );
  signal slice0_y_net_x3 : std_logic_vector( 16-1 downto 0 );
  signal slice1_y_net_x5 : std_logic_vector( 16-1 downto 0 );
  signal bitbasher4_a_net : std_logic_vector( 256-1 downto 0 );
  signal slice5_y_net_x2 : std_logic_vector( 16-1 downto 0 );
  signal slice5_y_net_x3 : std_logic_vector( 16-1 downto 0 );
  signal slice10_y_net_x4 : std_logic_vector( 16-1 downto 0 );
  signal slice3_y_net_x5 : std_logic_vector( 16-1 downto 0 );
  signal slice0_y_net_x5 : std_logic_vector( 16-1 downto 0 );
  signal slice15_y_net_x6 : std_logic_vector( 16-1 downto 0 );
  signal slice7_y_net_x4 : std_logic_vector( 16-1 downto 0 );
  signal slice14_y_net_x4 : std_logic_vector( 16-1 downto 0 );
  signal bitbasher3_a_net : std_logic_vector( 256-1 downto 0 );
  signal slice14_y_net_x5 : std_logic_vector( 16-1 downto 0 );
  signal slice13_y_net_x3 : std_logic_vector( 16-1 downto 0 );
  signal slice14_y_net_x3 : std_logic_vector( 16-1 downto 0 );
  signal slice12_y_net_x5 : std_logic_vector( 16-1 downto 0 );
  signal slice12_y_net_x4 : std_logic_vector( 16-1 downto 0 );
  signal slice4_y_net_x2 : std_logic_vector( 16-1 downto 0 );
  signal slice8_y_net_x1 : std_logic_vector( 16-1 downto 0 );
  signal slice8_y_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal slice12_y_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal slice0_y_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal slice0_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice8_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice3_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice10_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice15_y_net : std_logic_vector( 16-1 downto 0 );
  signal mux29_y_net : std_logic_vector( 17-1 downto 0 );
  signal mux37_y_net : std_logic_vector( 17-1 downto 0 );
  signal slice2_y_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal mux41_y_net : std_logic_vector( 17-1 downto 0 );
  signal slice9_y_net : std_logic_vector( 16-1 downto 0 );
  signal mux45_y_net : std_logic_vector( 17-1 downto 0 );
  signal slice0_y_net_x1 : std_logic_vector( 16-1 downto 0 );
  signal slice1_y_net_x1 : std_logic_vector( 16-1 downto 0 );
  signal slice10_y_net_x1 : std_logic_vector( 16-1 downto 0 );
  signal slice3_y_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal slice2_y_net_x1 : std_logic_vector( 16-1 downto 0 );
  signal slice10_y_net_x2 : std_logic_vector( 16-1 downto 0 );
  signal slice3_y_net_x1 : std_logic_vector( 16-1 downto 0 );
  signal slice14_y_net_x1 : std_logic_vector( 16-1 downto 0 );
  signal slice15_y_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal slice4_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice12_y_net_x2 : std_logic_vector( 16-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice1_y_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal slice5_y_net_x1 : std_logic_vector( 16-1 downto 0 );
  signal slice11_y_net_x1 : std_logic_vector( 16-1 downto 0 );
  signal slice13_y_net_x2 : std_logic_vector( 16-1 downto 0 );
  signal slice13_y_net_x1 : std_logic_vector( 16-1 downto 0 );
  signal slice13_y_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal slice5_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice7_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice15_y_net_x1 : std_logic_vector( 16-1 downto 0 );
  signal slice11_y_net_x2 : std_logic_vector( 16-1 downto 0 );
  signal bitbasher6_a_net : std_logic_vector( 256-1 downto 0 );
  signal slice14_y_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice4_y_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal slice6_y_net_x1 : std_logic_vector( 16-1 downto 0 );
  signal slice14_y_net_x2 : std_logic_vector( 16-1 downto 0 );
  signal slice11_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice13_y_net : std_logic_vector( 16-1 downto 0 );
  signal bitbasher7_a_net : std_logic_vector( 256-1 downto 0 );
  signal slice6_y_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal slice12_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice14_y_net : std_logic_vector( 16-1 downto 0 );
  signal bitbasher8_a_net : std_logic_vector( 256-1 downto 0 );
  signal slice6_y_net : std_logic_vector( 16-1 downto 0 );
  signal slice12_y_net_x1 : std_logic_vector( 16-1 downto 0 );
  signal mux2_y_net_x1 : std_logic_vector( 17-1 downto 0 );
  signal mux33_y_net : std_logic_vector( 17-1 downto 0 );
  signal slice7_y_net_x1 : std_logic_vector( 16-1 downto 0 );
  signal slice15_y_net_x2 : std_logic_vector( 16-1 downto 0 );
  signal slice9_y_net_x1 : std_logic_vector( 16-1 downto 0 );
  signal slice7_y_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal bitbasher5_a_net : std_logic_vector( 256-1 downto 0 );
  signal slice10_y_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal slice4_y_net_x1 : std_logic_vector( 16-1 downto 0 );
  signal slice5_y_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal slice9_y_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal slice11_y_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal constant7_op_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret16_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal reinterpret17_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal reinterpret19_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal reinterpret20_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal mux2_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret22_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal reinterpret1_output_port_net_x26 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net_x26 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net_x25 : std_logic_vector( 16-1 downto 0 );
  signal mux4_y_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal mux38_y_net : std_logic_vector( 17-1 downto 0 );
  signal mux30_y_net : std_logic_vector( 17-1 downto 0 );
  signal reinterpret29_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal constant3_op_net : std_logic_vector( 16-1 downto 0 );
  signal mux27_y_net : std_logic_vector( 17-1 downto 0 );
  signal mux50_y_net : std_logic_vector( 17-1 downto 0 );
  signal reinterpret25_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal reinterpret30_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 12-1 downto 0 );
  signal reinterpret26_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal reinterpret27_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal constant5_op_net : std_logic_vector( 16-1 downto 0 );
  signal mux7_y_net : std_logic_vector( 16-1 downto 0 );
  signal constant0_op_net : std_logic_vector( 16-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 12-1 downto 0 );
  signal reinterpret18_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 16-1 downto 0 );
  signal mux1_y_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal constant6_op_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret23_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal mux3_y_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal mux6_y_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal mux2_y_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal mux3_y_net : std_logic_vector( 16-1 downto 0 );
  signal mux5_y_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal mux4_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret21_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal delay9_q_net : std_logic_vector( 12-1 downto 0 );
  signal mux53_y_net : std_logic_vector( 17-1 downto 0 );
  signal delay10_q_net : std_logic_vector( 12-1 downto 0 );
  signal mux34_y_net : std_logic_vector( 17-1 downto 0 );
  signal delay11_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay12_q_net : std_logic_vector( 8-1 downto 0 );
  signal mux7_y_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal mux54_y_net : std_logic_vector( 17-1 downto 0 );
  signal mux49_y_net : std_logic_vector( 17-1 downto 0 );
  signal constant4_op_net : std_logic_vector( 16-1 downto 0 );
  signal delay16_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux0_y_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 16-1 downto 0 );
  signal mux5_y_net : std_logic_vector( 16-1 downto 0 );
  signal mux42_y_net : std_logic_vector( 17-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 12-1 downto 0 );
  signal reinterpret31_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal reinterpret24_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal delay11_q_net_x0 : std_logic_vector( 12-1 downto 0 );
  signal constant2_op_net : std_logic_vector( 16-1 downto 0 );
  signal mux46_y_net : std_logic_vector( 17-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 12-1 downto 0 );
  signal reinterpret28_output_port_net : std_logic_vector( 20-1 downto 0 );
  signal delay7_q_net : std_logic_vector( 12-1 downto 0 );
  signal mux0_y_net : std_logic_vector( 16-1 downto 0 );
  signal mux6_y_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net_x25 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net_x24 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net_x25 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net_x23 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net_x23 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net_x23 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net_x22 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net_x26 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net_x25 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net_x24 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net_x25 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net_x24 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net_x24 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net_x22 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net_x25 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net_x24 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net_x23 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net_x23 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net_x23 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net_x23 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net_x25 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net_x24 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net_x24 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net_x24 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net_x23 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net_x24 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net_x23 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net_x26 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net_x25 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net_x14 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net_x24 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net_x25 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net_x23 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net_x25 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net_x23 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net_x24 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net_x22 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net_x25 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net_x25 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net_x25 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net_x24 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net_x23 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net_x22 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net_x25 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net_x23 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net_x23 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net_x22 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net_x22 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net_x23 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net_x24 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net_x23 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net_x22 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net_x24 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net_x22 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net_x21 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net_x22 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net_x22 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net_x25 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net_x24 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net_x26 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net_x24 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net_x26 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net_x26 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net_x25 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net_x10 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net_x20 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net_x21 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net_x19 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net_x20 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net_x18 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net_x22 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net_x21 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net_x10 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net_x21 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net_x21 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net_x22 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net_x20 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net_x19 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net_x19 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net_x22 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net_x21 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net_x19 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net_x19 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net_x22 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net_x20 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net_x20 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net_x22 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net_x21 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net_x21 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net_x20 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net_x20 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net_x19 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net_x21 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net_x19 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net_x21 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net_x20 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net_x19 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net_x19 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net_x19 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net_x20 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net_x19 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net_x19 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net_x19 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net_x19 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net_x21 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net_x21 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net_x21 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net_x20 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net_x20 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net_x20 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net_x21 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net_x20 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net_x18 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net_x19 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net_x19 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net_x18 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net_x21 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net_x20 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net_x21 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net_x22 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net_x20 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net_x18 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net_x18 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net_x18 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net_x20 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net_x18 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net_x18 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net_x10 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net_x10 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net_x7 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net_x7 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net_x7 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net_x9 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net_x9 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net_x10 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net_x9 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net_x7 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net_x7 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net_x7 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net_x9 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net_x7 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net_x7 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net_x7 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net_x10 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net_x10 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net_x9 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net_x9 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net_x6 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net_x6 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net_x6 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net_x6 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net_x6 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net_x9 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net_x10 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net_x6 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net_x6 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net_x7 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net_x7 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net_x10 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net_x9 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net_x6 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net_x6 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net_x6 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net_x10 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net_x3 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net_x10 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net_x3 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net_x6 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net_x9 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net_x7 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net_x6 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net_x6 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net_x6 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net_x10 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net_x9 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net_x7 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net_x6 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net_x3 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net_x9 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net_x7 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net_x6 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net_x10 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net_x9 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net_x10 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net_x9 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net_x10 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net_x9 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net_x9 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net_x10 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net_x9 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net_x7 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net_x7 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net_x2 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net_x3 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net_x2 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net_x2 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal concat1_y_net_x6 : std_logic_vector( 256-1 downto 0 );
  signal reinterpret6_output_port_net_x2 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net_x3 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net_x2 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net_x2 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net_x2 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net_x3 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net_x2 : std_logic_vector( 16-1 downto 0 );
  signal concat1_y_net_x5 : std_logic_vector( 256-1 downto 0 );
  signal reinterpret6_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net_x3 : std_logic_vector( 16-1 downto 0 );
  signal concat1_y_net_x4 : std_logic_vector( 256-1 downto 0 );
  signal reinterpret7_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret12_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net_x3 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net_x3 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net_x3 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net_x2 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret0_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret4_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net_x3 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net_x3 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net_x3 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret1_output_port_net_x2 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net_x2 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret9_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret6_output_port_net_x3 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net_x3 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret14_output_port_net_x2 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret5_output_port_net_x2 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret7_output_port_net_x2 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret13_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret11_output_port_net_x0 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret15_output_port_net_x2 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal reinterpret8_output_port_net_x3 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret3_output_port_net_x2 : std_logic_vector( 16-1 downto 0 );
  signal reinterpret10_output_port_net : std_logic_vector( 16-1 downto 0 );
  signal constant15_op_net : std_logic_vector( 11-1 downto 0 );
  signal test_systolicfft_vhdl_black_box_vo_net : std_logic;
  signal delay19_q_net : std_logic_vector( 1-1 downto 0 );
  signal fifo4_dout_net : std_logic_vector( 256-1 downto 0 );
  signal bitbasher3_b_net : std_logic_vector( 16-1 downto 0 );
  signal fifo1_dout_net : std_logic_vector( 256-1 downto 0 );
  signal register_q_net_x8 : std_logic_vector( 1-1 downto 0 );
  signal concat1_y_net_x1 : std_logic_vector( 256-1 downto 0 );
  signal concat1_y_net_x0 : std_logic_vector( 256-1 downto 0 );
  signal register_q_net_x9 : std_logic_vector( 1-1 downto 0 );
  signal concat1_y_net_x3 : std_logic_vector( 256-1 downto 0 );
  signal fifo3_dout_net : std_logic_vector( 256-1 downto 0 );
  signal bitbasher4_b_net : std_logic_vector( 16-1 downto 0 );
  signal bitbasher6_b_net : std_logic_vector( 16-1 downto 0 );
  signal fifo2_dout_net : std_logic_vector( 256-1 downto 0 );
  signal fifo6_dout_net : std_logic_vector( 256-1 downto 0 );
  signal concat1_y_net : std_logic_vector( 256-1 downto 0 );
  signal concat1_y_net_x2 : std_logic_vector( 256-1 downto 0 );
  signal bitbasher2_b_net : std_logic_vector( 16-1 downto 0 );
  signal fifo7_dout_net : std_logic_vector( 256-1 downto 0 );
  signal bitbasher1_b_net : std_logic_vector( 16-1 downto 0 );
  signal bitbasher5_b_net : std_logic_vector( 16-1 downto 0 );
  signal constant14_op_net : std_logic_vector( 1-1 downto 0 );
  signal bitbasher8_b_net : std_logic_vector( 16-1 downto 0 );
  signal constant16_op_net : std_logic_vector( 1-1 downto 0 );
  signal fifo5_dout_net : std_logic_vector( 256-1 downto 0 );
  signal constant2_op_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal constant6_op_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal constant1_op_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal constant4_op_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal constant3_op_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal bitbasher7_b_net : std_logic_vector( 16-1 downto 0 );
  signal fifo8_dout_net : std_logic_vector( 256-1 downto 0 );
  signal constant5_op_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay18_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay17_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay13_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay15_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay28_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay29_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay30_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay55_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay56_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay53_q_net : std_logic_vector( 1-1 downto 0 );
  signal fifo1_full_net : std_logic;
  signal fifo1_empty_net : std_logic;
  signal fifo8_empty_net : std_logic;
  signal fifo8_full_net : std_logic;
  signal fifo7_full_net : std_logic;
  signal fifo7_empty_net : std_logic;
begin
  gin_tl_reset_net <= gin_tl_reset;
  gin_tl_start_net <= gin_tl_start;
  gin_addr_net <= gin_addr;
  gin_dphi_net <= gin_dphi;
  gin_init_im_net <= gin_init_im;
  gin_init_re_net <= gin_init_re;
  gin_we_even_1_net <= gin_we_even_1;
  gin_we_even_2_net <= gin_we_even_2;
  gin_we_even_3_net <= gin_we_even_3;
  gin_we_even_4_net <= gin_we_even_4;
  gin_we_odd_1_net <= gin_we_odd_1;
  gin_we_odd_2_net <= gin_we_odd_2;
  gin_we_odd_3_net <= gin_we_odd_3;
  gin_we_odd_4_net <= gin_we_odd_4;
  gout_cordic_delay_even_1 <= counter1_op_net_x6;
  gout_psb_tvalid <= delay54_q_net;
  gout_delay_ifft <= counter1_op_net_x7;
  gout_ov_ifft <= expression_dout_net;
  gout_ov_add <= expression1_dout_net;
  ts_0_net <= ts_0;
  ts_1_net <= ts_1;
  ts_2_net <= ts_2;
  ts_3_net <= ts_3;
  ts_4_net <= ts_4;
  ts_5_net <= ts_5;
  ts_6_net <= ts_6;
  ts_7_net <= ts_7;
  ts_a_net <= ts_a;
  ts_w_net <= ts_w;
  gout_psb_im_0 <= reinterpret3_output_port_net_x14;
  gout_psb_im_1 <= reinterpret2_output_port_net_x14;
  gout_psb_im_2 <= reinterpret7_output_port_net_x14;
  gout_psb_im_3 <= reinterpret6_output_port_net_x14;
  gout_psb_re_0 <= reinterpret_output_port_net;
  gout_psb_re_1 <= reinterpret1_output_port_net_x14;
  gout_psb_re_2 <= reinterpret4_output_port_net_x14;
  gout_psb_re_3 <= reinterpret5_output_port_net_x14;
  clk_net <= clk_1;
  ce_net <= ce_1;
  x0001 : entity xil_defaultlib.psb3_0_0001 
  port map (
    rst => gin_tl_reset_net,
    en => gin_tl_start_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    out_x0 => register_q_net_x7
  );
  baseband_even_1 : entity xil_defaultlib.psb3_0_baseband_even_1 
  port map (
    in_tvalid => delay14_q_net,
    addr_r => ram_dphi_addr_op_net,
    addr_w => delay38_q_net,
    init_im_even => delay44_q_net,
    init_re_even => delay35_q_net,
    dphi_even => delay37_q_net,
    we => delay1_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    delay_count => counter1_op_net_x6,
    out_im => cordic_6_0_even_1_m_axis_dout_tdata_imag_net_x0,
    out_re => cordic_6_0_even_1_m_axis_dout_tdata_real_net_x0,
    out_tvalid => cordic_6_0_even_1_m_axis_dout_tvalid_net_x0
  );
  baseband_even_2 : entity xil_defaultlib.psb3_0_baseband_even_2 
  port map (
    in_tvalid => delay14_q_net,
    addr_r => ram_dphi_addr_op_net,
    addr_w => delay38_q_net,
    init_im_even_2 => delay44_q_net,
    init_re_even_2 => delay35_q_net,
    dphi_even_2 => delay37_q_net,
    we => delay8_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    out_im => cordic_6_0_even_2_m_axis_dout_tdata_imag_net_x0,
    out_re => cordic_6_0_even_2_m_axis_dout_tdata_real_net_x0
  );
  baseband_even_3 : entity xil_defaultlib.psb3_0_baseband_even_3 
  port map (
    in_tvalid => delay14_q_net,
    addr_r => ram_dphi_addr_op_net,
    addr_w => delay38_q_net,
    init_im_even => delay44_q_net,
    init_re_even => delay35_q_net,
    dphi_even => delay37_q_net,
    we => delay31_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    out_im => cordic_6_0_even_1_m_axis_dout_tdata_imag_net,
    out_re => cordic_6_0_even_1_m_axis_dout_tdata_real_net
  );
  baseband_even_4 : entity xil_defaultlib.psb3_0_baseband_even_4 
  port map (
    in_tvalid => delay14_q_net,
    addr_r => ram_dphi_addr_op_net,
    addr_w => delay38_q_net,
    init_im_even_2 => delay44_q_net,
    init_re_even_2 => delay35_q_net,
    dphi_even_2 => delay37_q_net,
    we => delay49_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    out_im => cordic_6_0_even_2_m_axis_dout_tdata_imag_net,
    out_re => cordic_6_0_even_2_m_axis_dout_tdata_real_net
  );
  baseband_odd_1 : entity xil_defaultlib.psb3_0_baseband_odd_1 
  port map (
    tvalid => delay14_q_net,
    addr_r => ram_dphi_addr_op_net,
    addr_w => delay38_q_net,
    init_im_odd => delay44_q_net,
    init_re_odd => delay35_q_net,
    dphi_odd => delay37_q_net,
    we => delay6_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    out_im => cordic_6_0_odd_1_m_axis_dout_tdata_imag_net_x0,
    out_re => cordic_6_0_odd_1_m_axis_dout_tdata_real_net_x0
  );
  baseband_odd_2 : entity xil_defaultlib.psb3_0_baseband_odd_2 
  port map (
    tvalid => delay14_q_net,
    addr_r => ram_dphi_addr_op_net,
    addr_w => delay38_q_net,
    init_im_odd_2 => delay44_q_net,
    init_re_odd_2 => delay35_q_net,
    dphi_odd_2 => delay37_q_net,
    we => delay26_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    out_im => cordic_6_0_odd_2_m_axis_dout_tdata_imag_net_x0,
    out_re => cordic_6_0_odd_2_m_axis_dout_tdata_real_net_x0
  );
  baseband_odd_3 : entity xil_defaultlib.psb3_0_baseband_odd_3 
  port map (
    tvalid => delay14_q_net,
    addr_r => ram_dphi_addr_op_net,
    addr_w => delay38_q_net,
    init_im_odd => delay44_q_net,
    init_re_odd => delay35_q_net,
    dphi_odd => delay37_q_net,
    we => delay48_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    out_im => cordic_6_0_odd_1_m_axis_dout_tdata_imag_net,
    out_re => cordic_6_0_odd_1_m_axis_dout_tdata_real_net
  );
  baseband_odd_4 : entity xil_defaultlib.psb3_0_baseband_odd_4 
  port map (
    tvalid => delay14_q_net,
    addr_r => ram_dphi_addr_op_net,
    addr_w => delay38_q_net,
    init_im_odd_2 => delay44_q_net,
    init_re_odd_2 => delay35_q_net,
    dphi_odd_2 => delay37_q_net,
    we => delay43_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    out_im => cordic_6_0_odd_2_m_axis_dout_tdata_imag_net,
    out_re => cordic_6_0_odd_2_m_axis_dout_tdata_real_net
  );
  dpram_fir_coeffs_1 : entity xil_defaultlib.psb3_0_dpram_fir_coeffs_1 
  port map (
    in_rst => gin_tl_reset_net,
    in_en => delay8_q_net_x3,
    clk_1 => clk_net,
    ce_1 => ce_net,
    out_fir_coeffs_1 => reinterpret0_output_port_net_x17,
    out_fir_coeffs_2 => reinterpret1_output_port_net_x18,
    out_fir_coeffs_3 => reinterpret2_output_port_net_x18,
    out_fir_coeffs_4 => reinterpret3_output_port_net_x18,
    out_fir_coeffs_5 => reinterpret4_output_port_net_x18,
    out_fir_coeffs_6 => reinterpret5_output_port_net_x18,
    out_fir_coeffs_7 => reinterpret6_output_port_net_x18,
    out_fir_coeffs_8 => reinterpret7_output_port_net_x18,
    out_fir_coeffs_9 => reinterpret8_output_port_net_x18,
    out_fir_coeffs_10 => reinterpret9_output_port_net_x17,
    out_fir_coeffs_11 => reinterpret10_output_port_net_x17,
    out_fir_coeffs_12 => reinterpret11_output_port_net_x17,
    out_fir_coeffs_13 => reinterpret12_output_port_net_x17,
    out_fir_coeffs_14 => reinterpret13_output_port_net_x17,
    out_fir_coeffs_15 => reinterpret14_output_port_net_x17,
    out_fir_coeffs_16 => reinterpret15_output_port_net_x17
  );
  dpram_fir_coeffs_2 : entity xil_defaultlib.psb3_0_dpram_fir_coeffs_2 
  port map (
    in_rst => gin_tl_reset_net,
    in_en => delay8_q_net_x3,
    clk_1 => clk_net,
    ce_1 => ce_net,
    out_fir_coeffs_1 => reinterpret0_output_port_net_x16,
    out_fir_coeffs_2 => reinterpret1_output_port_net_x17,
    out_fir_coeffs_3 => reinterpret2_output_port_net_x17,
    out_fir_coeffs_4 => reinterpret3_output_port_net_x17,
    out_fir_coeffs_5 => reinterpret4_output_port_net_x17,
    out_fir_coeffs_6 => reinterpret5_output_port_net_x17,
    out_fir_coeffs_7 => reinterpret6_output_port_net_x17,
    out_fir_coeffs_8 => reinterpret7_output_port_net_x17,
    out_fir_coeffs_9 => reinterpret8_output_port_net_x17,
    out_fir_coeffs_10 => reinterpret9_output_port_net_x16,
    out_fir_coeffs_11 => reinterpret10_output_port_net_x16,
    out_fir_coeffs_12 => reinterpret11_output_port_net_x16,
    out_fir_coeffs_13 => reinterpret12_output_port_net_x16,
    out_fir_coeffs_14 => reinterpret13_output_port_net_x16,
    out_fir_coeffs_15 => reinterpret14_output_port_net_x16,
    out_fir_coeffs_16 => reinterpret15_output_port_net_x16
  );
  dpram_fir_coeffs_3 : entity xil_defaultlib.psb3_0_dpram_fir_coeffs_3 
  port map (
    in_rst => gin_tl_reset_net,
    in_en => delay8_q_net_x3,
    clk_1 => clk_net,
    ce_1 => ce_net,
    out_fir_coeffs_1 => reinterpret0_output_port_net_x15,
    out_fir_coeffs_2 => reinterpret1_output_port_net_x16,
    out_fir_coeffs_3 => reinterpret2_output_port_net_x16,
    out_fir_coeffs_4 => reinterpret3_output_port_net_x16,
    out_fir_coeffs_5 => reinterpret4_output_port_net_x16,
    out_fir_coeffs_6 => reinterpret5_output_port_net_x16,
    out_fir_coeffs_7 => reinterpret6_output_port_net_x16,
    out_fir_coeffs_8 => reinterpret7_output_port_net_x16,
    out_fir_coeffs_9 => reinterpret8_output_port_net_x16,
    out_fir_coeffs_10 => reinterpret9_output_port_net_x15,
    out_fir_coeffs_11 => reinterpret10_output_port_net_x15,
    out_fir_coeffs_12 => reinterpret11_output_port_net_x15,
    out_fir_coeffs_13 => reinterpret12_output_port_net_x15,
    out_fir_coeffs_14 => reinterpret13_output_port_net_x15,
    out_fir_coeffs_15 => reinterpret14_output_port_net_x15,
    out_fir_coeffs_16 => reinterpret15_output_port_net_x15
  );
  dpram_fir_coeffs_4 : entity xil_defaultlib.psb3_0_dpram_fir_coeffs_4 
  port map (
    in_rst => gin_tl_reset_net,
    in_en => delay8_q_net_x3,
    clk_1 => clk_net,
    ce_1 => ce_net,
    out_fir_coeffs_1 => reinterpret0_output_port_net_x14,
    out_fir_coeffs_2 => reinterpret1_output_port_net_x15,
    out_fir_coeffs_3 => reinterpret2_output_port_net_x15,
    out_fir_coeffs_4 => reinterpret3_output_port_net_x15,
    out_fir_coeffs_5 => reinterpret4_output_port_net_x15,
    out_fir_coeffs_6 => reinterpret5_output_port_net_x15,
    out_fir_coeffs_7 => reinterpret6_output_port_net_x15,
    out_fir_coeffs_8 => reinterpret7_output_port_net_x15,
    out_fir_coeffs_9 => reinterpret8_output_port_net_x15,
    out_fir_coeffs_10 => reinterpret9_output_port_net_x14,
    out_fir_coeffs_11 => reinterpret10_output_port_net_x14,
    out_fir_coeffs_12 => reinterpret11_output_port_net_x14,
    out_fir_coeffs_13 => reinterpret12_output_port_net_x14,
    out_fir_coeffs_14 => reinterpret13_output_port_net_x14,
    out_fir_coeffs_15 => reinterpret14_output_port_net_x14,
    out_fir_coeffs_16 => reinterpret15_output_port_net_x14
  );
  overflow_detector_add_im_1 : entity xil_defaultlib.psb3_0_overflow_detector_add_im_1 
  port map (
    rst => gin_tl_reset_net,
    a_1 => mult0_p_net_x6,
    b_1 => reinterpret0_output_port_net_x4,
    s_1 => addsub0_s_net_x5,
    a_2 => mult1_p_net_x6,
    a_3 => mult2_p_net_x6,
    a_4 => mult3_p_net_x6,
    a_5 => mult4_p_net_x6,
    a_6 => mult5_p_net_x6,
    a_7 => mult6_p_net_x6,
    a_8 => mult7_p_net_x6,
    a_9 => mult8_p_net_x6,
    a_10 => mult9_p_net_x6,
    a_11 => mult10_p_net_x6,
    a_12 => mult11_p_net_x6,
    a_13 => mult12_p_net_x6,
    a_14 => mult13_p_net_x6,
    a_15 => mult14_p_net_x6,
    a_16 => mult15_p_net_x6,
    b_2 => reinterpret1_output_port_net_x4,
    b_3 => reinterpret2_output_port_net_x4,
    b_4 => reinterpret3_output_port_net_x4,
    b_5 => reinterpret4_output_port_net_x4,
    b_6 => reinterpret5_output_port_net_x4,
    b_7 => reinterpret6_output_port_net_x4,
    b_8 => reinterpret7_output_port_net_x4,
    b_9 => reinterpret8_output_port_net_x4,
    b_10 => reinterpret9_output_port_net_x4,
    b_11 => reinterpret10_output_port_net_x4,
    b_12 => reinterpret11_output_port_net_x4,
    b_13 => reinterpret12_output_port_net_x4,
    b_14 => reinterpret13_output_port_net_x4,
    b_15 => reinterpret14_output_port_net_x4,
    b_16 => reinterpret15_output_port_net_x4,
    s_2 => addsub1_s_net_x5,
    s_3 => addsub2_s_net_x5,
    s_4 => addsub3_s_net_x5,
    s_5 => addsub4_s_net_x5,
    s_6 => addsub5_s_net_x5,
    s_7 => addsub6_s_net_x4,
    s_8 => addsub7_s_net_x5,
    s_9 => addsub8_s_net_x5,
    s_10 => addsub9_s_net_x5,
    s_11 => addsub10_s_net_x5,
    s_12 => addsub11_s_net_x5,
    s_13 => addsub12_s_net_x5,
    s_14 => addsub13_s_net_x5,
    s_15 => addsub14_s_net_x5,
    s_16 => addsub15_s_net_x5,
    clk_1 => clk_net,
    ce_1 => ce_net,
    ov => register_q_net_x6
  );
  overflow_detector_add_im_2 : entity xil_defaultlib.psb3_0_overflow_detector_add_im_2 
  port map (
    rst => gin_tl_reset_net,
    a_1 => mult0_p_net_x5,
    b_1 => reinterpret0_output_port_net_x1,
    s_1 => addsub0_s_net_x3,
    a_2 => mult1_p_net_x5,
    a_3 => mult2_p_net_x5,
    a_4 => mult3_p_net_x5,
    a_5 => mult4_p_net_x5,
    a_6 => mult5_p_net_x5,
    a_7 => mult6_p_net_x5,
    a_8 => mult7_p_net_x5,
    a_9 => mult8_p_net_x5,
    a_10 => mult9_p_net_x5,
    a_11 => mult10_p_net_x5,
    a_12 => mult11_p_net_x5,
    a_13 => mult12_p_net_x5,
    a_14 => mult13_p_net_x5,
    a_15 => mult14_p_net_x5,
    a_16 => mult15_p_net_x5,
    b_2 => reinterpret1_output_port_net_x1,
    b_3 => reinterpret2_output_port_net_x1,
    b_4 => reinterpret3_output_port_net_x1,
    b_5 => reinterpret4_output_port_net_x1,
    b_6 => reinterpret5_output_port_net_x1,
    b_7 => reinterpret6_output_port_net_x1,
    b_8 => reinterpret7_output_port_net_x1,
    b_9 => reinterpret8_output_port_net_x1,
    b_10 => reinterpret9_output_port_net_x1,
    b_11 => reinterpret10_output_port_net_x1,
    b_12 => reinterpret11_output_port_net_x1,
    b_13 => reinterpret12_output_port_net_x1,
    b_14 => reinterpret13_output_port_net_x1,
    b_15 => reinterpret14_output_port_net_x1,
    b_16 => reinterpret15_output_port_net_x1,
    s_2 => addsub1_s_net_x3,
    s_3 => addsub2_s_net_x3,
    s_4 => addsub3_s_net_x3,
    s_5 => addsub4_s_net_x3,
    s_6 => addsub5_s_net_x3,
    s_7 => addsub6_s_net_x2,
    s_8 => addsub7_s_net_x3,
    s_9 => addsub8_s_net_x3,
    s_10 => addsub9_s_net_x3,
    s_11 => addsub10_s_net_x3,
    s_12 => addsub11_s_net_x3,
    s_13 => addsub12_s_net_x3,
    s_14 => addsub13_s_net_x3,
    s_15 => addsub14_s_net_x3,
    s_16 => addsub15_s_net_x3,
    clk_1 => clk_net,
    ce_1 => ce_net,
    ov => register_q_net_x5
  );
  overflow_detector_add_im_3 : entity xil_defaultlib.psb3_0_overflow_detector_add_im_3 
  port map (
    rst => gin_tl_reset_net,
    a_1 => mult0_p_net_x4,
    b_1 => reinterpret0_output_port_net_x11,
    s_1 => addsub0_s_net_x1,
    a_2 => mult1_p_net_x4,
    a_3 => mult2_p_net_x4,
    a_4 => mult3_p_net_x4,
    a_5 => mult4_p_net_x4,
    a_6 => mult5_p_net_x4,
    a_7 => mult6_p_net_x4,
    a_8 => mult7_p_net_x4,
    a_9 => mult8_p_net_x4,
    a_10 => mult9_p_net_x4,
    a_11 => mult10_p_net_x4,
    a_12 => mult11_p_net_x4,
    a_13 => mult12_p_net_x4,
    a_14 => mult13_p_net_x4,
    a_15 => mult14_p_net_x4,
    a_16 => mult15_p_net_x4,
    b_2 => reinterpret1_output_port_net_x11,
    b_3 => reinterpret2_output_port_net_x11,
    b_4 => reinterpret3_output_port_net_x11,
    b_5 => reinterpret4_output_port_net_x11,
    b_6 => reinterpret5_output_port_net_x11,
    b_7 => reinterpret6_output_port_net_x11,
    b_8 => reinterpret7_output_port_net_x11,
    b_9 => reinterpret8_output_port_net_x11,
    b_10 => reinterpret9_output_port_net_x11,
    b_11 => reinterpret10_output_port_net_x11,
    b_12 => reinterpret11_output_port_net_x11,
    b_13 => reinterpret12_output_port_net_x11,
    b_14 => reinterpret13_output_port_net_x11,
    b_15 => reinterpret14_output_port_net_x11,
    b_16 => reinterpret15_output_port_net_x11,
    s_2 => addsub1_s_net_x1,
    s_3 => addsub2_s_net_x1,
    s_4 => addsub3_s_net_x1,
    s_5 => addsub4_s_net_x1,
    s_6 => addsub5_s_net_x1,
    s_7 => addsub6_s_net_x6,
    s_8 => addsub7_s_net_x1,
    s_9 => addsub8_s_net_x1,
    s_10 => addsub9_s_net_x1,
    s_11 => addsub10_s_net_x1,
    s_12 => addsub11_s_net_x1,
    s_13 => addsub12_s_net_x1,
    s_14 => addsub13_s_net_x1,
    s_15 => addsub14_s_net_x1,
    s_16 => addsub15_s_net_x1,
    clk_1 => clk_net,
    ce_1 => ce_net,
    ov => register_q_net_x4
  );
  overflow_detector_add_im_4 : entity xil_defaultlib.psb3_0_overflow_detector_add_im_4 
  port map (
    rst => gin_tl_reset_net,
    a_1 => mult0_p_net_x3,
    b_1 => reinterpret0_output_port_net_x8,
    s_1 => addsub0_s_net,
    a_2 => mult1_p_net_x3,
    a_3 => mult2_p_net_x3,
    a_4 => mult3_p_net_x3,
    a_5 => mult4_p_net_x3,
    a_6 => mult5_p_net_x3,
    a_7 => mult6_p_net_x3,
    a_8 => mult7_p_net_x3,
    a_9 => mult8_p_net_x3,
    a_10 => mult9_p_net_x3,
    a_11 => mult10_p_net_x3,
    a_12 => mult11_p_net_x3,
    a_13 => mult12_p_net_x3,
    a_14 => mult13_p_net_x3,
    a_15 => mult14_p_net_x3,
    a_16 => mult15_p_net_x3,
    b_2 => reinterpret1_output_port_net_x8,
    b_3 => reinterpret2_output_port_net_x8,
    b_4 => reinterpret3_output_port_net_x8,
    b_5 => reinterpret4_output_port_net_x8,
    b_6 => reinterpret5_output_port_net_x8,
    b_7 => reinterpret6_output_port_net_x8,
    b_8 => reinterpret7_output_port_net_x8,
    b_9 => reinterpret8_output_port_net_x8,
    b_10 => reinterpret9_output_port_net_x8,
    b_11 => reinterpret10_output_port_net_x8,
    b_12 => reinterpret11_output_port_net_x8,
    b_13 => reinterpret12_output_port_net_x8,
    b_14 => reinterpret13_output_port_net_x8,
    b_15 => reinterpret14_output_port_net_x8,
    b_16 => reinterpret15_output_port_net_x8,
    s_2 => addsub1_s_net,
    s_3 => addsub2_s_net,
    s_4 => addsub3_s_net,
    s_5 => addsub4_s_net,
    s_6 => addsub5_s_net,
    s_7 => addsub6_s_net,
    s_8 => addsub7_s_net,
    s_9 => addsub8_s_net,
    s_10 => addsub9_s_net,
    s_11 => addsub10_s_net,
    s_12 => addsub11_s_net,
    s_13 => addsub12_s_net,
    s_14 => addsub13_s_net,
    s_15 => addsub14_s_net,
    s_16 => addsub15_s_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    ov => register_q_net_x3
  );
  overflow_detector_add_re_1 : entity xil_defaultlib.psb3_0_overflow_detector_add_re_1 
  port map (
    rst => gin_tl_reset_net,
    a_1 => mult0_p_net_x2,
    b_1 => reinterpret0_output_port_net_x5,
    s_1 => addsub0_s_net_x6,
    a_2 => mult1_p_net_x2,
    a_3 => mult2_p_net_x2,
    a_4 => mult3_p_net_x2,
    a_5 => mult4_p_net_x2,
    a_6 => mult5_p_net_x2,
    a_7 => mult6_p_net_x2,
    a_8 => mult7_p_net_x2,
    a_9 => mult8_p_net_x2,
    a_10 => mult9_p_net_x2,
    a_11 => mult10_p_net_x2,
    a_12 => mult11_p_net_x2,
    a_13 => mult12_p_net_x2,
    a_14 => mult13_p_net_x2,
    a_15 => mult14_p_net_x2,
    a_16 => mult15_p_net_x2,
    b_2 => reinterpret1_output_port_net_x5,
    b_3 => reinterpret2_output_port_net_x5,
    b_4 => reinterpret3_output_port_net_x5,
    b_5 => reinterpret4_output_port_net_x5,
    b_6 => reinterpret5_output_port_net_x5,
    b_7 => reinterpret6_output_port_net_x5,
    b_8 => reinterpret7_output_port_net_x5,
    b_9 => reinterpret8_output_port_net_x5,
    b_10 => reinterpret9_output_port_net_x5,
    b_11 => reinterpret10_output_port_net_x5,
    b_12 => reinterpret11_output_port_net_x5,
    b_13 => reinterpret12_output_port_net_x5,
    b_14 => reinterpret13_output_port_net_x5,
    b_15 => reinterpret14_output_port_net_x5,
    b_16 => reinterpret15_output_port_net_x5,
    s_2 => addsub1_s_net_x6,
    s_3 => addsub2_s_net_x6,
    s_4 => addsub3_s_net_x6,
    s_5 => addsub4_s_net_x6,
    s_6 => addsub5_s_net_x6,
    s_7 => addsub6_s_net_x5,
    s_8 => addsub7_s_net_x6,
    s_9 => addsub8_s_net_x6,
    s_10 => addsub9_s_net_x6,
    s_11 => addsub10_s_net_x6,
    s_12 => addsub11_s_net_x6,
    s_13 => addsub12_s_net_x6,
    s_14 => addsub13_s_net_x6,
    s_15 => addsub14_s_net_x6,
    s_16 => addsub15_s_net_x6,
    clk_1 => clk_net,
    ce_1 => ce_net,
    ov => register_q_net_x2
  );
  overflow_detector_add_re_2 : entity xil_defaultlib.psb3_0_overflow_detector_add_re_2 
  port map (
    rst => gin_tl_reset_net,
    a_1 => mult0_p_net_x1,
    b_1 => reinterpret0_output_port_net_x13,
    s_1 => addsub0_s_net_x4,
    a_2 => mult1_p_net_x1,
    a_3 => mult2_p_net_x1,
    a_4 => mult3_p_net_x1,
    a_5 => mult4_p_net_x1,
    a_6 => mult5_p_net_x1,
    a_7 => mult6_p_net_x1,
    a_8 => mult7_p_net_x1,
    a_9 => mult8_p_net_x1,
    a_10 => mult9_p_net_x1,
    a_11 => mult10_p_net_x1,
    a_12 => mult11_p_net_x1,
    a_13 => mult12_p_net_x1,
    a_14 => mult13_p_net_x1,
    a_15 => mult14_p_net_x1,
    a_16 => mult15_p_net_x1,
    b_2 => reinterpret1_output_port_net_x13,
    b_3 => reinterpret2_output_port_net_x13,
    b_4 => reinterpret3_output_port_net_x13,
    b_5 => reinterpret4_output_port_net_x13,
    b_6 => reinterpret5_output_port_net_x13,
    b_7 => reinterpret6_output_port_net_x13,
    b_8 => reinterpret7_output_port_net_x13,
    b_9 => reinterpret8_output_port_net_x13,
    b_10 => reinterpret9_output_port_net_x13,
    b_11 => reinterpret10_output_port_net_x13,
    b_12 => reinterpret11_output_port_net_x13,
    b_13 => reinterpret12_output_port_net_x13,
    b_14 => reinterpret13_output_port_net_x13,
    b_15 => reinterpret14_output_port_net_x13,
    b_16 => reinterpret15_output_port_net_x13,
    s_2 => addsub1_s_net_x4,
    s_3 => addsub2_s_net_x4,
    s_4 => addsub3_s_net_x4,
    s_5 => addsub4_s_net_x4,
    s_6 => addsub5_s_net_x4,
    s_7 => addsub6_s_net_x3,
    s_8 => addsub7_s_net_x4,
    s_9 => addsub8_s_net_x4,
    s_10 => addsub9_s_net_x4,
    s_11 => addsub10_s_net_x4,
    s_12 => addsub11_s_net_x4,
    s_13 => addsub12_s_net_x4,
    s_14 => addsub13_s_net_x4,
    s_15 => addsub14_s_net_x4,
    s_16 => addsub15_s_net_x4,
    clk_1 => clk_net,
    ce_1 => ce_net,
    ov => register_q_net_x1
  );
  overflow_detector_add_re_3 : entity xil_defaultlib.psb3_0_overflow_detector_add_re_3 
  port map (
    rst => gin_tl_reset_net,
    a_1 => mult0_p_net_x0,
    b_1 => reinterpret0_output_port_net_x12,
    s_1 => addsub0_s_net_x2,
    a_2 => mult1_p_net_x0,
    a_3 => mult2_p_net_x0,
    a_4 => mult3_p_net_x0,
    a_5 => mult4_p_net_x0,
    a_6 => mult5_p_net_x0,
    a_7 => mult6_p_net_x0,
    a_8 => mult7_p_net_x0,
    a_9 => mult8_p_net_x0,
    a_10 => mult9_p_net_x0,
    a_11 => mult10_p_net_x0,
    a_12 => mult11_p_net_x0,
    a_13 => mult12_p_net_x0,
    a_14 => mult13_p_net_x0,
    a_15 => mult14_p_net_x0,
    a_16 => mult15_p_net_x0,
    b_2 => reinterpret1_output_port_net_x12,
    b_3 => reinterpret2_output_port_net_x12,
    b_4 => reinterpret3_output_port_net_x12,
    b_5 => reinterpret4_output_port_net_x12,
    b_6 => reinterpret5_output_port_net_x12,
    b_7 => reinterpret6_output_port_net_x12,
    b_8 => reinterpret7_output_port_net_x12,
    b_9 => reinterpret8_output_port_net_x12,
    b_10 => reinterpret9_output_port_net_x12,
    b_11 => reinterpret10_output_port_net_x12,
    b_12 => reinterpret11_output_port_net_x12,
    b_13 => reinterpret12_output_port_net_x12,
    b_14 => reinterpret13_output_port_net_x12,
    b_15 => reinterpret14_output_port_net_x12,
    b_16 => reinterpret15_output_port_net_x12,
    s_2 => addsub1_s_net_x2,
    s_3 => addsub2_s_net_x2,
    s_4 => addsub3_s_net_x2,
    s_5 => addsub4_s_net_x2,
    s_6 => addsub5_s_net_x2,
    s_7 => addsub6_s_net_x1,
    s_8 => addsub7_s_net_x2,
    s_9 => addsub8_s_net_x2,
    s_10 => addsub9_s_net_x2,
    s_11 => addsub10_s_net_x2,
    s_12 => addsub11_s_net_x2,
    s_13 => addsub12_s_net_x2,
    s_14 => addsub13_s_net_x2,
    s_15 => addsub14_s_net_x2,
    s_16 => addsub15_s_net_x2,
    clk_1 => clk_net,
    ce_1 => ce_net,
    ov => register_q_net_x0
  );
  overflow_detector_add_re_4 : entity xil_defaultlib.psb3_0_overflow_detector_add_re_4 
  port map (
    rst => gin_tl_reset_net,
    a_1 => mult0_p_net,
    b_1 => reinterpret0_output_port_net_x26,
    s_1 => addsub0_s_net_x0,
    a_2 => mult1_p_net,
    a_3 => mult2_p_net,
    a_4 => mult3_p_net,
    a_5 => mult4_p_net,
    a_6 => mult5_p_net,
    a_7 => mult6_p_net,
    a_8 => mult7_p_net,
    a_9 => mult8_p_net,
    a_10 => mult9_p_net,
    a_11 => mult10_p_net,
    a_12 => mult11_p_net,
    a_13 => mult12_p_net,
    a_14 => mult13_p_net,
    a_15 => mult14_p_net,
    a_16 => mult15_p_net,
    b_2 => reinterpret1_output_port_net_x27,
    b_3 => reinterpret2_output_port_net_x27,
    b_4 => reinterpret3_output_port_net_x27,
    b_5 => reinterpret4_output_port_net_x27,
    b_6 => reinterpret5_output_port_net_x27,
    b_7 => reinterpret6_output_port_net_x27,
    b_8 => reinterpret7_output_port_net_x27,
    b_9 => reinterpret8_output_port_net_x26,
    b_10 => reinterpret9_output_port_net_x26,
    b_11 => reinterpret10_output_port_net_x26,
    b_12 => reinterpret11_output_port_net_x26,
    b_13 => reinterpret12_output_port_net_x26,
    b_14 => reinterpret13_output_port_net_x26,
    b_15 => reinterpret14_output_port_net_x26,
    b_16 => reinterpret15_output_port_net_x26,
    s_2 => addsub1_s_net_x0,
    s_3 => addsub2_s_net_x0,
    s_4 => addsub3_s_net_x0,
    s_5 => addsub4_s_net_x0,
    s_6 => addsub5_s_net_x0,
    s_7 => addsub6_s_net_x0,
    s_8 => addsub7_s_net_x0,
    s_9 => addsub8_s_net_x0,
    s_10 => addsub9_s_net_x0,
    s_11 => addsub10_s_net_x0,
    s_12 => addsub11_s_net_x0,
    s_13 => addsub12_s_net_x0,
    s_14 => addsub13_s_net_x0,
    s_15 => addsub14_s_net_x0,
    s_16 => addsub15_s_net_x0,
    clk_1 => clk_net,
    ce_1 => ce_net,
    ov => register_q_net
  );
  scalar_to_vector1 : entity xil_defaultlib.psb3_0_scalar_to_vector1 
  port map (
    i => bitbasher1_a_net,
    o_1 => slice0_y_net_x6,
    o_2 => slice1_y_net_x6,
    o_3 => slice2_y_net_x6,
    o_4 => slice3_y_net_x6,
    o_5 => slice4_y_net_x6,
    o_6 => slice5_y_net_x6,
    o_7 => slice6_y_net_x6,
    o_8 => slice7_y_net_x6,
    o_9 => slice8_y_net_x6,
    o_10 => slice9_y_net_x6,
    o_11 => slice10_y_net_x6,
    o_12 => slice11_y_net_x6,
    o_13 => slice12_y_net_x6,
    o_14 => slice13_y_net_x6,
    o_15 => slice14_y_net_x6,
    o_16 => slice15_y_net_x6
  );
  scalar_to_vector2 : entity xil_defaultlib.psb3_0_scalar_to_vector2 
  port map (
    i => bitbasher2_a_net,
    o_1 => slice0_y_net_x5,
    o_2 => slice1_y_net_x5,
    o_3 => slice2_y_net_x5,
    o_4 => slice3_y_net_x5,
    o_5 => slice4_y_net_x5,
    o_6 => slice5_y_net_x5,
    o_7 => slice6_y_net_x5,
    o_8 => slice7_y_net_x5,
    o_9 => slice8_y_net_x5,
    o_10 => slice9_y_net_x5,
    o_11 => slice10_y_net_x5,
    o_12 => slice11_y_net_x5,
    o_13 => slice12_y_net_x5,
    o_14 => slice13_y_net_x5,
    o_15 => slice14_y_net_x5,
    o_16 => slice15_y_net_x5
  );
  scalar_to_vector3 : entity xil_defaultlib.psb3_0_scalar_to_vector3 
  port map (
    i => bitbasher3_a_net,
    o_1 => slice0_y_net_x4,
    o_2 => slice1_y_net_x4,
    o_3 => slice2_y_net_x4,
    o_4 => slice3_y_net_x4,
    o_5 => slice4_y_net_x4,
    o_6 => slice5_y_net_x4,
    o_7 => slice6_y_net_x4,
    o_8 => slice7_y_net_x4,
    o_9 => slice8_y_net_x4,
    o_10 => slice9_y_net_x4,
    o_11 => slice10_y_net_x4,
    o_12 => slice11_y_net_x4,
    o_13 => slice12_y_net_x4,
    o_14 => slice13_y_net_x4,
    o_15 => slice14_y_net_x4,
    o_16 => slice15_y_net_x4
  );
  scalar_to_vector4 : entity xil_defaultlib.psb3_0_scalar_to_vector4 
  port map (
    i => bitbasher4_a_net,
    o_1 => slice0_y_net_x3,
    o_2 => slice1_y_net_x3,
    o_3 => slice2_y_net_x3,
    o_4 => slice3_y_net_x3,
    o_5 => slice4_y_net_x3,
    o_6 => slice5_y_net_x3,
    o_7 => slice6_y_net_x3,
    o_8 => slice7_y_net_x3,
    o_9 => slice8_y_net_x3,
    o_10 => slice9_y_net_x3,
    o_11 => slice10_y_net_x3,
    o_12 => slice11_y_net_x3,
    o_13 => slice12_y_net_x3,
    o_14 => slice13_y_net_x3,
    o_15 => slice14_y_net_x3,
    o_16 => slice15_y_net_x3
  );
  scalar_to_vector5 : entity xil_defaultlib.psb3_0_scalar_to_vector5 
  port map (
    i => bitbasher5_a_net,
    o_1 => slice0_y_net_x2,
    o_2 => slice1_y_net_x2,
    o_3 => slice2_y_net_x2,
    o_4 => slice3_y_net_x2,
    o_5 => slice4_y_net_x2,
    o_6 => slice5_y_net_x2,
    o_7 => slice6_y_net_x2,
    o_8 => slice7_y_net_x2,
    o_9 => slice8_y_net_x2,
    o_10 => slice9_y_net_x2,
    o_11 => slice10_y_net_x2,
    o_12 => slice11_y_net_x2,
    o_13 => slice12_y_net_x2,
    o_14 => slice13_y_net_x2,
    o_15 => slice14_y_net_x2,
    o_16 => slice15_y_net_x2
  );
  scalar_to_vector6 : entity xil_defaultlib.psb3_0_scalar_to_vector6 
  port map (
    i => bitbasher6_a_net,
    o_1 => slice0_y_net_x1,
    o_2 => slice1_y_net_x1,
    o_3 => slice2_y_net_x1,
    o_4 => slice3_y_net_x1,
    o_5 => slice4_y_net_x1,
    o_6 => slice5_y_net_x1,
    o_7 => slice6_y_net_x1,
    o_8 => slice7_y_net_x1,
    o_9 => slice8_y_net_x1,
    o_10 => slice9_y_net_x1,
    o_11 => slice10_y_net_x1,
    o_12 => slice11_y_net_x1,
    o_13 => slice12_y_net_x1,
    o_14 => slice13_y_net_x1,
    o_15 => slice14_y_net_x1,
    o_16 => slice15_y_net_x1
  );
  scalar_to_vector7 : entity xil_defaultlib.psb3_0_scalar_to_vector7 
  port map (
    i => bitbasher7_a_net,
    o_1 => slice0_y_net_x0,
    o_2 => slice1_y_net_x0,
    o_3 => slice2_y_net_x0,
    o_4 => slice3_y_net_x0,
    o_5 => slice4_y_net_x0,
    o_6 => slice5_y_net_x0,
    o_7 => slice6_y_net_x0,
    o_8 => slice7_y_net_x0,
    o_9 => slice8_y_net_x0,
    o_10 => slice9_y_net_x0,
    o_11 => slice10_y_net_x0,
    o_12 => slice11_y_net_x0,
    o_13 => slice12_y_net_x0,
    o_14 => slice13_y_net_x0,
    o_15 => slice14_y_net_x0,
    o_16 => slice15_y_net_x0
  );
  scalar_to_vector8 : entity xil_defaultlib.psb3_0_scalar_to_vector8 
  port map (
    i => bitbasher8_a_net,
    o_1 => slice0_y_net,
    o_2 => slice1_y_net,
    o_3 => slice2_y_net,
    o_4 => slice3_y_net,
    o_5 => slice4_y_net,
    o_6 => slice5_y_net,
    o_7 => slice6_y_net,
    o_8 => slice7_y_net,
    o_9 => slice8_y_net,
    o_10 => slice9_y_net,
    o_11 => slice10_y_net,
    o_12 => slice11_y_net,
    o_13 => slice12_y_net,
    o_14 => slice13_y_net,
    o_15 => slice14_y_net,
    o_16 => slice15_y_net
  );
  toneselect : entity xil_defaultlib.psb3_0_toneselect 
  port map (
    in_even1_im => cordic_6_0_even_1_m_axis_dout_tdata_imag_net_x0,
    in_even1_re => cordic_6_0_even_1_m_axis_dout_tdata_real_net_x0,
    in_odd1_im => cordic_6_0_odd_1_m_axis_dout_tdata_imag_net_x0,
    in_odd1_re => cordic_6_0_odd_1_m_axis_dout_tdata_real_net_x0,
    in_even2_im => cordic_6_0_even_2_m_axis_dout_tdata_imag_net_x0,
    in_even2_re => cordic_6_0_even_2_m_axis_dout_tdata_real_net_x0,
    in_odd2_im => cordic_6_0_odd_2_m_axis_dout_tdata_imag_net_x0,
    in_odd2_re => cordic_6_0_odd_2_m_axis_dout_tdata_real_net_x0,
    in_even3_im => cordic_6_0_even_1_m_axis_dout_tdata_imag_net,
    in_even3_re => cordic_6_0_even_1_m_axis_dout_tdata_real_net,
    in_odd3_im => cordic_6_0_odd_1_m_axis_dout_tdata_imag_net,
    in_odd3_re => cordic_6_0_odd_1_m_axis_dout_tdata_real_net,
    in_even4_im => cordic_6_0_even_2_m_axis_dout_tdata_imag_net,
    in_even4_re => cordic_6_0_even_2_m_axis_dout_tdata_real_net,
    in_odd4_im => cordic_6_0_odd_2_m_axis_dout_tdata_imag_net,
    in_odd4_re => cordic_6_0_odd_2_m_axis_dout_tdata_real_net,
    in_tvalid => cordic_6_0_even_1_m_axis_dout_tvalid_net_x0,
    rst => gin_tl_reset_net,
    data_0 => delay2_q_net,
    data_1 => delay3_q_net,
    data_2 => delay4_q_net,
    data_3 => delay5_q_net,
    data_4 => delay7_q_net,
    data_5 => delay9_q_net,
    data_6 => delay10_q_net,
    data_7 => delay11_q_net_x0,
    w_addr_x0 => delay12_q_net,
    we => delay16_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    out_even1_re => mux2_y_net_x1,
    out_odd1_re => mux29_y_net,
    out_even2_re => mux33_y_net,
    out_odd2_re => mux37_y_net,
    out_even3_re => mux41_y_net,
    out_odd3_re => mux45_y_net,
    out_even4_re => mux49_y_net,
    out_odd4_re => mux53_y_net,
    out_even1_im => mux27_y_net,
    out_odd1_im => mux30_y_net,
    out_even2_im => mux34_y_net,
    out_odd2_im => mux38_y_net,
    out_even3_im => mux42_y_net,
    out_odd3_im => mux46_y_net,
    out_even4_im => mux50_y_net,
    out_odd4_im => mux54_y_net,
    out_tvalid => delay11_q_net
  );
  vector_addsub_fabric : entity xil_defaultlib.psb3_0_vector_addsub_fabric 
  port map (
    a_1 => mult0_p_net_x2,
    b_1 => reinterpret0_output_port_net_x5,
    a_2 => mult1_p_net_x2,
    a_3 => mult2_p_net_x2,
    a_4 => mult3_p_net_x2,
    a_5 => mult4_p_net_x2,
    a_6 => mult5_p_net_x2,
    a_7 => mult6_p_net_x2,
    a_8 => mult7_p_net_x2,
    a_9 => mult8_p_net_x2,
    a_10 => mult9_p_net_x2,
    a_11 => mult10_p_net_x2,
    a_12 => mult11_p_net_x2,
    a_13 => mult12_p_net_x2,
    a_14 => mult13_p_net_x2,
    a_15 => mult14_p_net_x2,
    a_16 => mult15_p_net_x2,
    b_2 => reinterpret1_output_port_net_x5,
    b_3 => reinterpret2_output_port_net_x5,
    b_4 => reinterpret3_output_port_net_x5,
    b_5 => reinterpret4_output_port_net_x5,
    b_6 => reinterpret5_output_port_net_x5,
    b_7 => reinterpret6_output_port_net_x5,
    b_8 => reinterpret7_output_port_net_x5,
    b_9 => reinterpret8_output_port_net_x5,
    b_10 => reinterpret9_output_port_net_x5,
    b_11 => reinterpret10_output_port_net_x5,
    b_12 => reinterpret11_output_port_net_x5,
    b_13 => reinterpret12_output_port_net_x5,
    b_14 => reinterpret13_output_port_net_x5,
    b_15 => reinterpret14_output_port_net_x5,
    b_16 => reinterpret15_output_port_net_x5,
    clk_1 => clk_net,
    ce_1 => ce_net,
    a_b_1 => addsub0_s_net_x6,
    a_b_2 => addsub1_s_net_x6,
    a_b_3 => addsub2_s_net_x6,
    a_b_4 => addsub3_s_net_x6,
    a_b_5 => addsub4_s_net_x6,
    a_b_6 => addsub5_s_net_x6,
    a_b_7 => addsub6_s_net_x5,
    a_b_8 => addsub7_s_net_x6,
    a_b_9 => addsub8_s_net_x6,
    a_b_10 => addsub9_s_net_x6,
    a_b_11 => addsub10_s_net_x6,
    a_b_12 => addsub11_s_net_x6,
    a_b_13 => addsub12_s_net_x6,
    a_b_14 => addsub13_s_net_x6,
    a_b_15 => addsub14_s_net_x6,
    a_b_16 => addsub15_s_net_x6
  );
  vector_addsub_fabric1 : entity xil_defaultlib.psb3_0_vector_addsub_fabric1 
  port map (
    a_1 => mult0_p_net_x6,
    b_1 => reinterpret0_output_port_net_x4,
    a_2 => mult1_p_net_x6,
    a_3 => mult2_p_net_x6,
    a_4 => mult3_p_net_x6,
    a_5 => mult4_p_net_x6,
    a_6 => mult5_p_net_x6,
    a_7 => mult6_p_net_x6,
    a_8 => mult7_p_net_x6,
    a_9 => mult8_p_net_x6,
    a_10 => mult9_p_net_x6,
    a_11 => mult10_p_net_x6,
    a_12 => mult11_p_net_x6,
    a_13 => mult12_p_net_x6,
    a_14 => mult13_p_net_x6,
    a_15 => mult14_p_net_x6,
    a_16 => mult15_p_net_x6,
    b_2 => reinterpret1_output_port_net_x4,
    b_3 => reinterpret2_output_port_net_x4,
    b_4 => reinterpret3_output_port_net_x4,
    b_5 => reinterpret4_output_port_net_x4,
    b_6 => reinterpret5_output_port_net_x4,
    b_7 => reinterpret6_output_port_net_x4,
    b_8 => reinterpret7_output_port_net_x4,
    b_9 => reinterpret8_output_port_net_x4,
    b_10 => reinterpret9_output_port_net_x4,
    b_11 => reinterpret10_output_port_net_x4,
    b_12 => reinterpret11_output_port_net_x4,
    b_13 => reinterpret12_output_port_net_x4,
    b_14 => reinterpret13_output_port_net_x4,
    b_15 => reinterpret14_output_port_net_x4,
    b_16 => reinterpret15_output_port_net_x4,
    clk_1 => clk_net,
    ce_1 => ce_net,
    a_b_1 => addsub0_s_net_x5,
    a_b_2 => addsub1_s_net_x5,
    a_b_3 => addsub2_s_net_x5,
    a_b_4 => addsub3_s_net_x5,
    a_b_5 => addsub4_s_net_x5,
    a_b_6 => addsub5_s_net_x5,
    a_b_7 => addsub6_s_net_x4,
    a_b_8 => addsub7_s_net_x5,
    a_b_9 => addsub8_s_net_x5,
    a_b_10 => addsub9_s_net_x5,
    a_b_11 => addsub10_s_net_x5,
    a_b_12 => addsub11_s_net_x5,
    a_b_13 => addsub12_s_net_x5,
    a_b_14 => addsub13_s_net_x5,
    a_b_15 => addsub14_s_net_x5,
    a_b_16 => addsub15_s_net_x5
  );
  vector_addsub_fabric2 : entity xil_defaultlib.psb3_0_vector_addsub_fabric2 
  port map (
    a_1 => mult0_p_net_x1,
    b_1 => reinterpret0_output_port_net_x13,
    a_2 => mult1_p_net_x1,
    a_3 => mult2_p_net_x1,
    a_4 => mult3_p_net_x1,
    a_5 => mult4_p_net_x1,
    a_6 => mult5_p_net_x1,
    a_7 => mult6_p_net_x1,
    a_8 => mult7_p_net_x1,
    a_9 => mult8_p_net_x1,
    a_10 => mult9_p_net_x1,
    a_11 => mult10_p_net_x1,
    a_12 => mult11_p_net_x1,
    a_13 => mult12_p_net_x1,
    a_14 => mult13_p_net_x1,
    a_15 => mult14_p_net_x1,
    a_16 => mult15_p_net_x1,
    b_2 => reinterpret1_output_port_net_x13,
    b_3 => reinterpret2_output_port_net_x13,
    b_4 => reinterpret3_output_port_net_x13,
    b_5 => reinterpret4_output_port_net_x13,
    b_6 => reinterpret5_output_port_net_x13,
    b_7 => reinterpret6_output_port_net_x13,
    b_8 => reinterpret7_output_port_net_x13,
    b_9 => reinterpret8_output_port_net_x13,
    b_10 => reinterpret9_output_port_net_x13,
    b_11 => reinterpret10_output_port_net_x13,
    b_12 => reinterpret11_output_port_net_x13,
    b_13 => reinterpret12_output_port_net_x13,
    b_14 => reinterpret13_output_port_net_x13,
    b_15 => reinterpret14_output_port_net_x13,
    b_16 => reinterpret15_output_port_net_x13,
    clk_1 => clk_net,
    ce_1 => ce_net,
    a_b_1 => addsub0_s_net_x4,
    a_b_2 => addsub1_s_net_x4,
    a_b_3 => addsub2_s_net_x4,
    a_b_4 => addsub3_s_net_x4,
    a_b_5 => addsub4_s_net_x4,
    a_b_6 => addsub5_s_net_x4,
    a_b_7 => addsub6_s_net_x3,
    a_b_8 => addsub7_s_net_x4,
    a_b_9 => addsub8_s_net_x4,
    a_b_10 => addsub9_s_net_x4,
    a_b_11 => addsub10_s_net_x4,
    a_b_12 => addsub11_s_net_x4,
    a_b_13 => addsub12_s_net_x4,
    a_b_14 => addsub13_s_net_x4,
    a_b_15 => addsub14_s_net_x4,
    a_b_16 => addsub15_s_net_x4
  );
  vector_addsub_fabric3 : entity xil_defaultlib.psb3_0_vector_addsub_fabric3 
  port map (
    a_1 => mult0_p_net_x5,
    b_1 => reinterpret0_output_port_net_x1,
    a_2 => mult1_p_net_x5,
    a_3 => mult2_p_net_x5,
    a_4 => mult3_p_net_x5,
    a_5 => mult4_p_net_x5,
    a_6 => mult5_p_net_x5,
    a_7 => mult6_p_net_x5,
    a_8 => mult7_p_net_x5,
    a_9 => mult8_p_net_x5,
    a_10 => mult9_p_net_x5,
    a_11 => mult10_p_net_x5,
    a_12 => mult11_p_net_x5,
    a_13 => mult12_p_net_x5,
    a_14 => mult13_p_net_x5,
    a_15 => mult14_p_net_x5,
    a_16 => mult15_p_net_x5,
    b_2 => reinterpret1_output_port_net_x1,
    b_3 => reinterpret2_output_port_net_x1,
    b_4 => reinterpret3_output_port_net_x1,
    b_5 => reinterpret4_output_port_net_x1,
    b_6 => reinterpret5_output_port_net_x1,
    b_7 => reinterpret6_output_port_net_x1,
    b_8 => reinterpret7_output_port_net_x1,
    b_9 => reinterpret8_output_port_net_x1,
    b_10 => reinterpret9_output_port_net_x1,
    b_11 => reinterpret10_output_port_net_x1,
    b_12 => reinterpret11_output_port_net_x1,
    b_13 => reinterpret12_output_port_net_x1,
    b_14 => reinterpret13_output_port_net_x1,
    b_15 => reinterpret14_output_port_net_x1,
    b_16 => reinterpret15_output_port_net_x1,
    clk_1 => clk_net,
    ce_1 => ce_net,
    a_b_1 => addsub0_s_net_x3,
    a_b_2 => addsub1_s_net_x3,
    a_b_3 => addsub2_s_net_x3,
    a_b_4 => addsub3_s_net_x3,
    a_b_5 => addsub4_s_net_x3,
    a_b_6 => addsub5_s_net_x3,
    a_b_7 => addsub6_s_net_x2,
    a_b_8 => addsub7_s_net_x3,
    a_b_9 => addsub8_s_net_x3,
    a_b_10 => addsub9_s_net_x3,
    a_b_11 => addsub10_s_net_x3,
    a_b_12 => addsub11_s_net_x3,
    a_b_13 => addsub12_s_net_x3,
    a_b_14 => addsub13_s_net_x3,
    a_b_15 => addsub14_s_net_x3,
    a_b_16 => addsub15_s_net_x3
  );
  vector_addsub_fabric4 : entity xil_defaultlib.psb3_0_vector_addsub_fabric4 
  port map (
    a_1 => mult0_p_net_x0,
    b_1 => reinterpret0_output_port_net_x12,
    a_2 => mult1_p_net_x0,
    a_3 => mult2_p_net_x0,
    a_4 => mult3_p_net_x0,
    a_5 => mult4_p_net_x0,
    a_6 => mult5_p_net_x0,
    a_7 => mult6_p_net_x0,
    a_8 => mult7_p_net_x0,
    a_9 => mult8_p_net_x0,
    a_10 => mult9_p_net_x0,
    a_11 => mult10_p_net_x0,
    a_12 => mult11_p_net_x0,
    a_13 => mult12_p_net_x0,
    a_14 => mult13_p_net_x0,
    a_15 => mult14_p_net_x0,
    a_16 => mult15_p_net_x0,
    b_2 => reinterpret1_output_port_net_x12,
    b_3 => reinterpret2_output_port_net_x12,
    b_4 => reinterpret3_output_port_net_x12,
    b_5 => reinterpret4_output_port_net_x12,
    b_6 => reinterpret5_output_port_net_x12,
    b_7 => reinterpret6_output_port_net_x12,
    b_8 => reinterpret7_output_port_net_x12,
    b_9 => reinterpret8_output_port_net_x12,
    b_10 => reinterpret9_output_port_net_x12,
    b_11 => reinterpret10_output_port_net_x12,
    b_12 => reinterpret11_output_port_net_x12,
    b_13 => reinterpret12_output_port_net_x12,
    b_14 => reinterpret13_output_port_net_x12,
    b_15 => reinterpret14_output_port_net_x12,
    b_16 => reinterpret15_output_port_net_x12,
    clk_1 => clk_net,
    ce_1 => ce_net,
    a_b_1 => addsub0_s_net_x2,
    a_b_2 => addsub1_s_net_x2,
    a_b_3 => addsub2_s_net_x2,
    a_b_4 => addsub3_s_net_x2,
    a_b_5 => addsub4_s_net_x2,
    a_b_6 => addsub5_s_net_x2,
    a_b_7 => addsub6_s_net_x1,
    a_b_8 => addsub7_s_net_x2,
    a_b_9 => addsub8_s_net_x2,
    a_b_10 => addsub9_s_net_x2,
    a_b_11 => addsub10_s_net_x2,
    a_b_12 => addsub11_s_net_x2,
    a_b_13 => addsub12_s_net_x2,
    a_b_14 => addsub13_s_net_x2,
    a_b_15 => addsub14_s_net_x2,
    a_b_16 => addsub15_s_net_x2
  );
  vector_addsub_fabric5 : entity xil_defaultlib.psb3_0_vector_addsub_fabric5 
  port map (
    a_1 => mult0_p_net_x4,
    b_1 => reinterpret0_output_port_net_x11,
    a_2 => mult1_p_net_x4,
    a_3 => mult2_p_net_x4,
    a_4 => mult3_p_net_x4,
    a_5 => mult4_p_net_x4,
    a_6 => mult5_p_net_x4,
    a_7 => mult6_p_net_x4,
    a_8 => mult7_p_net_x4,
    a_9 => mult8_p_net_x4,
    a_10 => mult9_p_net_x4,
    a_11 => mult10_p_net_x4,
    a_12 => mult11_p_net_x4,
    a_13 => mult12_p_net_x4,
    a_14 => mult13_p_net_x4,
    a_15 => mult14_p_net_x4,
    a_16 => mult15_p_net_x4,
    b_2 => reinterpret1_output_port_net_x11,
    b_3 => reinterpret2_output_port_net_x11,
    b_4 => reinterpret3_output_port_net_x11,
    b_5 => reinterpret4_output_port_net_x11,
    b_6 => reinterpret5_output_port_net_x11,
    b_7 => reinterpret6_output_port_net_x11,
    b_8 => reinterpret7_output_port_net_x11,
    b_9 => reinterpret8_output_port_net_x11,
    b_10 => reinterpret9_output_port_net_x11,
    b_11 => reinterpret10_output_port_net_x11,
    b_12 => reinterpret11_output_port_net_x11,
    b_13 => reinterpret12_output_port_net_x11,
    b_14 => reinterpret13_output_port_net_x11,
    b_15 => reinterpret14_output_port_net_x11,
    b_16 => reinterpret15_output_port_net_x11,
    clk_1 => clk_net,
    ce_1 => ce_net,
    a_b_1 => addsub0_s_net_x1,
    a_b_2 => addsub1_s_net_x1,
    a_b_3 => addsub2_s_net_x1,
    a_b_4 => addsub3_s_net_x1,
    a_b_5 => addsub4_s_net_x1,
    a_b_6 => addsub5_s_net_x1,
    a_b_7 => addsub6_s_net_x6,
    a_b_8 => addsub7_s_net_x1,
    a_b_9 => addsub8_s_net_x1,
    a_b_10 => addsub9_s_net_x1,
    a_b_11 => addsub10_s_net_x1,
    a_b_12 => addsub11_s_net_x1,
    a_b_13 => addsub12_s_net_x1,
    a_b_14 => addsub13_s_net_x1,
    a_b_15 => addsub14_s_net_x1,
    a_b_16 => addsub15_s_net_x1
  );
  vector_addsub_fabric6 : entity xil_defaultlib.psb3_0_vector_addsub_fabric6 
  port map (
    a_1 => mult0_p_net,
    b_1 => reinterpret0_output_port_net_x26,
    a_2 => mult1_p_net,
    a_3 => mult2_p_net,
    a_4 => mult3_p_net,
    a_5 => mult4_p_net,
    a_6 => mult5_p_net,
    a_7 => mult6_p_net,
    a_8 => mult7_p_net,
    a_9 => mult8_p_net,
    a_10 => mult9_p_net,
    a_11 => mult10_p_net,
    a_12 => mult11_p_net,
    a_13 => mult12_p_net,
    a_14 => mult13_p_net,
    a_15 => mult14_p_net,
    a_16 => mult15_p_net,
    b_2 => reinterpret1_output_port_net_x27,
    b_3 => reinterpret2_output_port_net_x27,
    b_4 => reinterpret3_output_port_net_x27,
    b_5 => reinterpret4_output_port_net_x27,
    b_6 => reinterpret5_output_port_net_x27,
    b_7 => reinterpret6_output_port_net_x27,
    b_8 => reinterpret7_output_port_net_x27,
    b_9 => reinterpret8_output_port_net_x26,
    b_10 => reinterpret9_output_port_net_x26,
    b_11 => reinterpret10_output_port_net_x26,
    b_12 => reinterpret11_output_port_net_x26,
    b_13 => reinterpret12_output_port_net_x26,
    b_14 => reinterpret13_output_port_net_x26,
    b_15 => reinterpret14_output_port_net_x26,
    b_16 => reinterpret15_output_port_net_x26,
    clk_1 => clk_net,
    ce_1 => ce_net,
    a_b_1 => addsub0_s_net_x0,
    a_b_2 => addsub1_s_net_x0,
    a_b_3 => addsub2_s_net_x0,
    a_b_4 => addsub3_s_net_x0,
    a_b_5 => addsub4_s_net_x0,
    a_b_6 => addsub5_s_net_x0,
    a_b_7 => addsub6_s_net_x0,
    a_b_8 => addsub7_s_net_x0,
    a_b_9 => addsub8_s_net_x0,
    a_b_10 => addsub9_s_net_x0,
    a_b_11 => addsub10_s_net_x0,
    a_b_12 => addsub11_s_net_x0,
    a_b_13 => addsub12_s_net_x0,
    a_b_14 => addsub13_s_net_x0,
    a_b_15 => addsub14_s_net_x0,
    a_b_16 => addsub15_s_net_x0
  );
  vector_addsub_fabric7 : entity xil_defaultlib.psb3_0_vector_addsub_fabric7 
  port map (
    a_1 => mult0_p_net_x3,
    b_1 => reinterpret0_output_port_net_x8,
    a_2 => mult1_p_net_x3,
    a_3 => mult2_p_net_x3,
    a_4 => mult3_p_net_x3,
    a_5 => mult4_p_net_x3,
    a_6 => mult5_p_net_x3,
    a_7 => mult6_p_net_x3,
    a_8 => mult7_p_net_x3,
    a_9 => mult8_p_net_x3,
    a_10 => mult9_p_net_x3,
    a_11 => mult10_p_net_x3,
    a_12 => mult11_p_net_x3,
    a_13 => mult12_p_net_x3,
    a_14 => mult13_p_net_x3,
    a_15 => mult14_p_net_x3,
    a_16 => mult15_p_net_x3,
    b_2 => reinterpret1_output_port_net_x8,
    b_3 => reinterpret2_output_port_net_x8,
    b_4 => reinterpret3_output_port_net_x8,
    b_5 => reinterpret4_output_port_net_x8,
    b_6 => reinterpret5_output_port_net_x8,
    b_7 => reinterpret6_output_port_net_x8,
    b_8 => reinterpret7_output_port_net_x8,
    b_9 => reinterpret8_output_port_net_x8,
    b_10 => reinterpret9_output_port_net_x8,
    b_11 => reinterpret10_output_port_net_x8,
    b_12 => reinterpret11_output_port_net_x8,
    b_13 => reinterpret12_output_port_net_x8,
    b_14 => reinterpret13_output_port_net_x8,
    b_15 => reinterpret14_output_port_net_x8,
    b_16 => reinterpret15_output_port_net_x8,
    clk_1 => clk_net,
    ce_1 => ce_net,
    a_b_1 => addsub0_s_net,
    a_b_2 => addsub1_s_net,
    a_b_3 => addsub2_s_net,
    a_b_4 => addsub3_s_net,
    a_b_5 => addsub4_s_net,
    a_b_6 => addsub5_s_net,
    a_b_7 => addsub6_s_net,
    a_b_8 => addsub7_s_net,
    a_b_9 => addsub8_s_net,
    a_b_10 => addsub9_s_net,
    a_b_11 => addsub10_s_net,
    a_b_12 => addsub11_s_net,
    a_b_13 => addsub12_s_net,
    a_b_14 => addsub13_s_net,
    a_b_15 => addsub14_s_net,
    a_b_16 => addsub15_s_net
  );
  vector_constant : entity xil_defaultlib.psb3_0_vector_constant 
  port map (
    out1_1 => constant0_op_net,
    out1_2 => constant1_op_net,
    out1_3 => constant2_op_net,
    out1_4 => constant3_op_net,
    out1_5 => constant4_op_net,
    out1_6 => constant5_op_net,
    out1_7 => constant6_op_net,
    out1_8 => constant7_op_net
  );
  vector_mux : entity xil_defaultlib.psb3_0_vector_mux 
  port map (
    sel => register_q_net_x7,
    i0_1 => constant0_op_net,
    i1_1 => reinterpret24_output_port_net,
    i0_2 => constant1_op_net,
    i0_3 => constant2_op_net,
    i0_4 => constant3_op_net,
    i0_5 => constant4_op_net,
    i0_6 => constant5_op_net,
    i0_7 => constant6_op_net,
    i0_8 => constant7_op_net,
    i1_2 => reinterpret25_output_port_net,
    i1_3 => reinterpret26_output_port_net,
    i1_4 => reinterpret27_output_port_net,
    i1_5 => reinterpret28_output_port_net,
    i1_6 => reinterpret29_output_port_net,
    i1_7 => reinterpret30_output_port_net,
    i1_8 => reinterpret31_output_port_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    o_1 => mux0_y_net_x0,
    o_2 => mux1_y_net_x0,
    o_3 => mux2_y_net_x0,
    o_4 => mux3_y_net_x0,
    o_5 => mux4_y_net_x0,
    o_6 => mux5_y_net_x0,
    o_7 => mux6_y_net_x0,
    o_8 => mux7_y_net_x0
  );
  vector_mux1 : entity xil_defaultlib.psb3_0_vector_mux1 
  port map (
    sel => register_q_net_x7,
    i0_1 => constant0_op_net,
    i1_1 => reinterpret16_output_port_net,
    i0_2 => constant1_op_net,
    i0_3 => constant2_op_net,
    i0_4 => constant3_op_net,
    i0_5 => constant4_op_net,
    i0_6 => constant5_op_net,
    i0_7 => constant6_op_net,
    i0_8 => constant7_op_net,
    i1_2 => reinterpret17_output_port_net,
    i1_3 => reinterpret18_output_port_net,
    i1_4 => reinterpret19_output_port_net,
    i1_5 => reinterpret20_output_port_net,
    i1_6 => reinterpret21_output_port_net,
    i1_7 => reinterpret22_output_port_net,
    i1_8 => reinterpret23_output_port_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    o_1 => mux0_y_net,
    o_2 => mux1_y_net,
    o_3 => mux2_y_net,
    o_4 => mux3_y_net,
    o_5 => mux4_y_net,
    o_6 => mux5_y_net,
    o_7 => mux6_y_net,
    o_8 => mux7_y_net
  );
  vector_real_mult_im_1 : entity xil_defaultlib.psb3_0_vector_real_mult_im_1 
  port map (
    a_1 => reinterpret0_output_port_net_x25,
    b_1 => reinterpret0_output_port_net_x17,
    a_2 => reinterpret1_output_port_net_x26,
    a_3 => reinterpret2_output_port_net_x26,
    a_4 => reinterpret3_output_port_net_x26,
    a_5 => reinterpret4_output_port_net_x26,
    a_6 => reinterpret5_output_port_net_x26,
    a_7 => reinterpret6_output_port_net_x26,
    a_8 => reinterpret7_output_port_net_x26,
    a_9 => reinterpret8_output_port_net_x25,
    a_10 => reinterpret9_output_port_net_x25,
    a_11 => reinterpret10_output_port_net_x25,
    a_12 => reinterpret11_output_port_net_x25,
    a_13 => reinterpret12_output_port_net_x25,
    a_14 => reinterpret13_output_port_net_x25,
    a_15 => reinterpret14_output_port_net_x25,
    a_16 => reinterpret15_output_port_net_x25,
    b_2 => reinterpret1_output_port_net_x18,
    b_3 => reinterpret2_output_port_net_x18,
    b_4 => reinterpret3_output_port_net_x18,
    b_5 => reinterpret4_output_port_net_x18,
    b_6 => reinterpret5_output_port_net_x18,
    b_7 => reinterpret6_output_port_net_x18,
    b_8 => reinterpret7_output_port_net_x18,
    b_9 => reinterpret8_output_port_net_x18,
    b_10 => reinterpret9_output_port_net_x17,
    b_11 => reinterpret10_output_port_net_x17,
    b_12 => reinterpret11_output_port_net_x17,
    b_13 => reinterpret12_output_port_net_x17,
    b_14 => reinterpret13_output_port_net_x17,
    b_15 => reinterpret14_output_port_net_x17,
    b_16 => reinterpret15_output_port_net_x17,
    clk_1 => clk_net,
    ce_1 => ce_net,
    a_x_b_1 => mult0_p_net_x6,
    a_x_b_2 => mult1_p_net_x6,
    a_x_b_3 => mult2_p_net_x6,
    a_x_b_4 => mult3_p_net_x6,
    a_x_b_5 => mult4_p_net_x6,
    a_x_b_6 => mult5_p_net_x6,
    a_x_b_7 => mult6_p_net_x6,
    a_x_b_8 => mult7_p_net_x6,
    a_x_b_9 => mult8_p_net_x6,
    a_x_b_10 => mult9_p_net_x6,
    a_x_b_11 => mult10_p_net_x6,
    a_x_b_12 => mult11_p_net_x6,
    a_x_b_13 => mult12_p_net_x6,
    a_x_b_14 => mult13_p_net_x6,
    a_x_b_15 => mult14_p_net_x6,
    a_x_b_16 => mult15_p_net_x6
  );
  vector_real_mult_im_2 : entity xil_defaultlib.psb3_0_vector_real_mult_im_2 
  port map (
    a_1 => reinterpret0_output_port_net_x24,
    b_1 => reinterpret0_output_port_net_x16,
    a_2 => reinterpret1_output_port_net_x25,
    a_3 => reinterpret2_output_port_net_x25,
    a_4 => reinterpret3_output_port_net_x25,
    a_5 => reinterpret4_output_port_net_x25,
    a_6 => reinterpret5_output_port_net_x25,
    a_7 => reinterpret6_output_port_net_x25,
    a_8 => reinterpret7_output_port_net_x25,
    a_9 => reinterpret8_output_port_net_x14,
    a_10 => reinterpret9_output_port_net_x24,
    a_11 => reinterpret10_output_port_net_x24,
    a_12 => reinterpret11_output_port_net_x24,
    a_13 => reinterpret12_output_port_net_x24,
    a_14 => reinterpret13_output_port_net_x24,
    a_15 => reinterpret14_output_port_net_x24,
    a_16 => reinterpret15_output_port_net_x24,
    b_2 => reinterpret1_output_port_net_x17,
    b_3 => reinterpret2_output_port_net_x17,
    b_4 => reinterpret3_output_port_net_x17,
    b_5 => reinterpret4_output_port_net_x17,
    b_6 => reinterpret5_output_port_net_x17,
    b_7 => reinterpret6_output_port_net_x17,
    b_8 => reinterpret7_output_port_net_x17,
    b_9 => reinterpret8_output_port_net_x17,
    b_10 => reinterpret9_output_port_net_x16,
    b_11 => reinterpret10_output_port_net_x16,
    b_12 => reinterpret11_output_port_net_x16,
    b_13 => reinterpret12_output_port_net_x16,
    b_14 => reinterpret13_output_port_net_x16,
    b_15 => reinterpret14_output_port_net_x16,
    b_16 => reinterpret15_output_port_net_x16,
    clk_1 => clk_net,
    ce_1 => ce_net,
    a_x_b_1 => mult0_p_net_x5,
    a_x_b_2 => mult1_p_net_x5,
    a_x_b_3 => mult2_p_net_x5,
    a_x_b_4 => mult3_p_net_x5,
    a_x_b_5 => mult4_p_net_x5,
    a_x_b_6 => mult5_p_net_x5,
    a_x_b_7 => mult6_p_net_x5,
    a_x_b_8 => mult7_p_net_x5,
    a_x_b_9 => mult8_p_net_x5,
    a_x_b_10 => mult9_p_net_x5,
    a_x_b_11 => mult10_p_net_x5,
    a_x_b_12 => mult11_p_net_x5,
    a_x_b_13 => mult12_p_net_x5,
    a_x_b_14 => mult13_p_net_x5,
    a_x_b_15 => mult14_p_net_x5,
    a_x_b_16 => mult15_p_net_x5
  );
  vector_real_mult_im_3 : entity xil_defaultlib.psb3_0_vector_real_mult_im_3 
  port map (
    a_1 => reinterpret0_output_port_net_x23,
    b_1 => reinterpret0_output_port_net_x15,
    a_2 => reinterpret1_output_port_net_x24,
    a_3 => reinterpret2_output_port_net_x24,
    a_4 => reinterpret3_output_port_net_x24,
    a_5 => reinterpret4_output_port_net_x24,
    a_6 => reinterpret5_output_port_net_x24,
    a_7 => reinterpret6_output_port_net_x24,
    a_8 => reinterpret7_output_port_net_x24,
    a_9 => reinterpret8_output_port_net_x24,
    a_10 => reinterpret9_output_port_net_x23,
    a_11 => reinterpret10_output_port_net_x23,
    a_12 => reinterpret11_output_port_net_x23,
    a_13 => reinterpret12_output_port_net_x23,
    a_14 => reinterpret13_output_port_net_x23,
    a_15 => reinterpret14_output_port_net_x23,
    a_16 => reinterpret15_output_port_net_x23,
    b_2 => reinterpret1_output_port_net_x16,
    b_3 => reinterpret2_output_port_net_x16,
    b_4 => reinterpret3_output_port_net_x16,
    b_5 => reinterpret4_output_port_net_x16,
    b_6 => reinterpret5_output_port_net_x16,
    b_7 => reinterpret6_output_port_net_x16,
    b_8 => reinterpret7_output_port_net_x16,
    b_9 => reinterpret8_output_port_net_x16,
    b_10 => reinterpret9_output_port_net_x15,
    b_11 => reinterpret10_output_port_net_x15,
    b_12 => reinterpret11_output_port_net_x15,
    b_13 => reinterpret12_output_port_net_x15,
    b_14 => reinterpret13_output_port_net_x15,
    b_15 => reinterpret14_output_port_net_x15,
    b_16 => reinterpret15_output_port_net_x15,
    clk_1 => clk_net,
    ce_1 => ce_net,
    a_x_b_1 => mult0_p_net_x4,
    a_x_b_2 => mult1_p_net_x4,
    a_x_b_3 => mult2_p_net_x4,
    a_x_b_4 => mult3_p_net_x4,
    a_x_b_5 => mult4_p_net_x4,
    a_x_b_6 => mult5_p_net_x4,
    a_x_b_7 => mult6_p_net_x4,
    a_x_b_8 => mult7_p_net_x4,
    a_x_b_9 => mult8_p_net_x4,
    a_x_b_10 => mult9_p_net_x4,
    a_x_b_11 => mult10_p_net_x4,
    a_x_b_12 => mult11_p_net_x4,
    a_x_b_13 => mult12_p_net_x4,
    a_x_b_14 => mult13_p_net_x4,
    a_x_b_15 => mult14_p_net_x4,
    a_x_b_16 => mult15_p_net_x4
  );
  vector_real_mult_im_4 : entity xil_defaultlib.psb3_0_vector_real_mult_im_4 
  port map (
    a_1 => reinterpret0_output_port_net_x22,
    b_1 => reinterpret0_output_port_net_x14,
    a_2 => reinterpret1_output_port_net_x23,
    a_3 => reinterpret2_output_port_net_x23,
    a_4 => reinterpret3_output_port_net_x23,
    a_5 => reinterpret4_output_port_net_x23,
    a_6 => reinterpret5_output_port_net_x23,
    a_7 => reinterpret6_output_port_net_x23,
    a_8 => reinterpret7_output_port_net_x23,
    a_9 => reinterpret8_output_port_net_x23,
    a_10 => reinterpret9_output_port_net_x22,
    a_11 => reinterpret10_output_port_net_x22,
    a_12 => reinterpret11_output_port_net_x22,
    a_13 => reinterpret12_output_port_net_x22,
    a_14 => reinterpret13_output_port_net_x22,
    a_15 => reinterpret14_output_port_net_x22,
    a_16 => reinterpret15_output_port_net_x22,
    b_2 => reinterpret1_output_port_net_x15,
    b_3 => reinterpret2_output_port_net_x15,
    b_4 => reinterpret3_output_port_net_x15,
    b_5 => reinterpret4_output_port_net_x15,
    b_6 => reinterpret5_output_port_net_x15,
    b_7 => reinterpret6_output_port_net_x15,
    b_8 => reinterpret7_output_port_net_x15,
    b_9 => reinterpret8_output_port_net_x15,
    b_10 => reinterpret9_output_port_net_x14,
    b_11 => reinterpret10_output_port_net_x14,
    b_12 => reinterpret11_output_port_net_x14,
    b_13 => reinterpret12_output_port_net_x14,
    b_14 => reinterpret13_output_port_net_x14,
    b_15 => reinterpret14_output_port_net_x14,
    b_16 => reinterpret15_output_port_net_x14,
    clk_1 => clk_net,
    ce_1 => ce_net,
    a_x_b_1 => mult0_p_net_x3,
    a_x_b_2 => mult1_p_net_x3,
    a_x_b_3 => mult2_p_net_x3,
    a_x_b_4 => mult3_p_net_x3,
    a_x_b_5 => mult4_p_net_x3,
    a_x_b_6 => mult5_p_net_x3,
    a_x_b_7 => mult6_p_net_x3,
    a_x_b_8 => mult7_p_net_x3,
    a_x_b_9 => mult8_p_net_x3,
    a_x_b_10 => mult9_p_net_x3,
    a_x_b_11 => mult10_p_net_x3,
    a_x_b_12 => mult11_p_net_x3,
    a_x_b_13 => mult12_p_net_x3,
    a_x_b_14 => mult13_p_net_x3,
    a_x_b_15 => mult14_p_net_x3,
    a_x_b_16 => mult15_p_net_x3
  );
  vector_real_mult_re_1 : entity xil_defaultlib.psb3_0_vector_real_mult_re_1 
  port map (
    a_1 => reinterpret0_output_port_net_x21,
    b_1 => reinterpret0_output_port_net_x17,
    a_2 => reinterpret1_output_port_net_x22,
    a_3 => reinterpret2_output_port_net_x22,
    a_4 => reinterpret3_output_port_net_x22,
    a_5 => reinterpret4_output_port_net_x22,
    a_6 => reinterpret5_output_port_net_x22,
    a_7 => reinterpret6_output_port_net_x22,
    a_8 => reinterpret7_output_port_net_x22,
    a_9 => reinterpret8_output_port_net_x22,
    a_10 => reinterpret9_output_port_net_x21,
    a_11 => reinterpret10_output_port_net_x21,
    a_12 => reinterpret11_output_port_net_x21,
    a_13 => reinterpret12_output_port_net_x21,
    a_14 => reinterpret13_output_port_net_x21,
    a_15 => reinterpret14_output_port_net_x21,
    a_16 => reinterpret15_output_port_net_x21,
    b_2 => reinterpret1_output_port_net_x18,
    b_3 => reinterpret2_output_port_net_x18,
    b_4 => reinterpret3_output_port_net_x18,
    b_5 => reinterpret4_output_port_net_x18,
    b_6 => reinterpret5_output_port_net_x18,
    b_7 => reinterpret6_output_port_net_x18,
    b_8 => reinterpret7_output_port_net_x18,
    b_9 => reinterpret8_output_port_net_x18,
    b_10 => reinterpret9_output_port_net_x17,
    b_11 => reinterpret10_output_port_net_x17,
    b_12 => reinterpret11_output_port_net_x17,
    b_13 => reinterpret12_output_port_net_x17,
    b_14 => reinterpret13_output_port_net_x17,
    b_15 => reinterpret14_output_port_net_x17,
    b_16 => reinterpret15_output_port_net_x17,
    clk_1 => clk_net,
    ce_1 => ce_net,
    a_x_b_1 => mult0_p_net_x2,
    a_x_b_2 => mult1_p_net_x2,
    a_x_b_3 => mult2_p_net_x2,
    a_x_b_4 => mult3_p_net_x2,
    a_x_b_5 => mult4_p_net_x2,
    a_x_b_6 => mult5_p_net_x2,
    a_x_b_7 => mult6_p_net_x2,
    a_x_b_8 => mult7_p_net_x2,
    a_x_b_9 => mult8_p_net_x2,
    a_x_b_10 => mult9_p_net_x2,
    a_x_b_11 => mult10_p_net_x2,
    a_x_b_12 => mult11_p_net_x2,
    a_x_b_13 => mult12_p_net_x2,
    a_x_b_14 => mult13_p_net_x2,
    a_x_b_15 => mult14_p_net_x2,
    a_x_b_16 => mult15_p_net_x2
  );
  vector_real_mult_re_2 : entity xil_defaultlib.psb3_0_vector_real_mult_re_2 
  port map (
    a_1 => reinterpret0_output_port_net_x20,
    b_1 => reinterpret0_output_port_net_x16,
    a_2 => reinterpret1_output_port_net_x21,
    a_3 => reinterpret2_output_port_net_x21,
    a_4 => reinterpret3_output_port_net_x21,
    a_5 => reinterpret4_output_port_net_x21,
    a_6 => reinterpret5_output_port_net_x21,
    a_7 => reinterpret6_output_port_net_x21,
    a_8 => reinterpret7_output_port_net_x21,
    a_9 => reinterpret8_output_port_net_x21,
    a_10 => reinterpret9_output_port_net_x20,
    a_11 => reinterpret10_output_port_net_x20,
    a_12 => reinterpret11_output_port_net_x20,
    a_13 => reinterpret12_output_port_net_x20,
    a_14 => reinterpret13_output_port_net_x20,
    a_15 => reinterpret14_output_port_net_x20,
    a_16 => reinterpret15_output_port_net_x20,
    b_2 => reinterpret1_output_port_net_x17,
    b_3 => reinterpret2_output_port_net_x17,
    b_4 => reinterpret3_output_port_net_x17,
    b_5 => reinterpret4_output_port_net_x17,
    b_6 => reinterpret5_output_port_net_x17,
    b_7 => reinterpret6_output_port_net_x17,
    b_8 => reinterpret7_output_port_net_x17,
    b_9 => reinterpret8_output_port_net_x17,
    b_10 => reinterpret9_output_port_net_x16,
    b_11 => reinterpret10_output_port_net_x16,
    b_12 => reinterpret11_output_port_net_x16,
    b_13 => reinterpret12_output_port_net_x16,
    b_14 => reinterpret13_output_port_net_x16,
    b_15 => reinterpret14_output_port_net_x16,
    b_16 => reinterpret15_output_port_net_x16,
    clk_1 => clk_net,
    ce_1 => ce_net,
    a_x_b_1 => mult0_p_net_x1,
    a_x_b_2 => mult1_p_net_x1,
    a_x_b_3 => mult2_p_net_x1,
    a_x_b_4 => mult3_p_net_x1,
    a_x_b_5 => mult4_p_net_x1,
    a_x_b_6 => mult5_p_net_x1,
    a_x_b_7 => mult6_p_net_x1,
    a_x_b_8 => mult7_p_net_x1,
    a_x_b_9 => mult8_p_net_x1,
    a_x_b_10 => mult9_p_net_x1,
    a_x_b_11 => mult10_p_net_x1,
    a_x_b_12 => mult11_p_net_x1,
    a_x_b_13 => mult12_p_net_x1,
    a_x_b_14 => mult13_p_net_x1,
    a_x_b_15 => mult14_p_net_x1,
    a_x_b_16 => mult15_p_net_x1
  );
  vector_real_mult_re_3 : entity xil_defaultlib.psb3_0_vector_real_mult_re_3 
  port map (
    a_1 => reinterpret0_output_port_net_x19,
    b_1 => reinterpret0_output_port_net_x15,
    a_2 => reinterpret1_output_port_net_x20,
    a_3 => reinterpret2_output_port_net_x20,
    a_4 => reinterpret3_output_port_net_x20,
    a_5 => reinterpret4_output_port_net_x20,
    a_6 => reinterpret5_output_port_net_x20,
    a_7 => reinterpret6_output_port_net_x20,
    a_8 => reinterpret7_output_port_net_x20,
    a_9 => reinterpret8_output_port_net_x20,
    a_10 => reinterpret9_output_port_net_x19,
    a_11 => reinterpret10_output_port_net_x19,
    a_12 => reinterpret11_output_port_net_x19,
    a_13 => reinterpret12_output_port_net_x19,
    a_14 => reinterpret13_output_port_net_x19,
    a_15 => reinterpret14_output_port_net_x19,
    a_16 => reinterpret15_output_port_net_x19,
    b_2 => reinterpret1_output_port_net_x16,
    b_3 => reinterpret2_output_port_net_x16,
    b_4 => reinterpret3_output_port_net_x16,
    b_5 => reinterpret4_output_port_net_x16,
    b_6 => reinterpret5_output_port_net_x16,
    b_7 => reinterpret6_output_port_net_x16,
    b_8 => reinterpret7_output_port_net_x16,
    b_9 => reinterpret8_output_port_net_x16,
    b_10 => reinterpret9_output_port_net_x15,
    b_11 => reinterpret10_output_port_net_x15,
    b_12 => reinterpret11_output_port_net_x15,
    b_13 => reinterpret12_output_port_net_x15,
    b_14 => reinterpret13_output_port_net_x15,
    b_15 => reinterpret14_output_port_net_x15,
    b_16 => reinterpret15_output_port_net_x15,
    clk_1 => clk_net,
    ce_1 => ce_net,
    a_x_b_1 => mult0_p_net_x0,
    a_x_b_2 => mult1_p_net_x0,
    a_x_b_3 => mult2_p_net_x0,
    a_x_b_4 => mult3_p_net_x0,
    a_x_b_5 => mult4_p_net_x0,
    a_x_b_6 => mult5_p_net_x0,
    a_x_b_7 => mult6_p_net_x0,
    a_x_b_8 => mult7_p_net_x0,
    a_x_b_9 => mult8_p_net_x0,
    a_x_b_10 => mult9_p_net_x0,
    a_x_b_11 => mult10_p_net_x0,
    a_x_b_12 => mult11_p_net_x0,
    a_x_b_13 => mult12_p_net_x0,
    a_x_b_14 => mult13_p_net_x0,
    a_x_b_15 => mult14_p_net_x0,
    a_x_b_16 => mult15_p_net_x0
  );
  vector_real_mult_re_4 : entity xil_defaultlib.psb3_0_vector_real_mult_re_4 
  port map (
    a_1 => reinterpret0_output_port_net_x18,
    b_1 => reinterpret0_output_port_net_x14,
    a_2 => reinterpret1_output_port_net_x19,
    a_3 => reinterpret2_output_port_net_x19,
    a_4 => reinterpret3_output_port_net_x19,
    a_5 => reinterpret4_output_port_net_x19,
    a_6 => reinterpret5_output_port_net_x19,
    a_7 => reinterpret6_output_port_net_x19,
    a_8 => reinterpret7_output_port_net_x19,
    a_9 => reinterpret8_output_port_net_x19,
    a_10 => reinterpret9_output_port_net_x18,
    a_11 => reinterpret10_output_port_net_x18,
    a_12 => reinterpret11_output_port_net_x18,
    a_13 => reinterpret12_output_port_net_x18,
    a_14 => reinterpret13_output_port_net_x18,
    a_15 => reinterpret14_output_port_net_x18,
    a_16 => reinterpret15_output_port_net_x18,
    b_2 => reinterpret1_output_port_net_x15,
    b_3 => reinterpret2_output_port_net_x15,
    b_4 => reinterpret3_output_port_net_x15,
    b_5 => reinterpret4_output_port_net_x15,
    b_6 => reinterpret5_output_port_net_x15,
    b_7 => reinterpret6_output_port_net_x15,
    b_8 => reinterpret7_output_port_net_x15,
    b_9 => reinterpret8_output_port_net_x15,
    b_10 => reinterpret9_output_port_net_x14,
    b_11 => reinterpret10_output_port_net_x14,
    b_12 => reinterpret11_output_port_net_x14,
    b_13 => reinterpret12_output_port_net_x14,
    b_14 => reinterpret13_output_port_net_x14,
    b_15 => reinterpret14_output_port_net_x14,
    b_16 => reinterpret15_output_port_net_x14,
    clk_1 => clk_net,
    ce_1 => ce_net,
    a_x_b_1 => mult0_p_net,
    a_x_b_2 => mult1_p_net,
    a_x_b_3 => mult2_p_net,
    a_x_b_4 => mult3_p_net,
    a_x_b_5 => mult4_p_net,
    a_x_b_6 => mult5_p_net,
    a_x_b_7 => mult6_p_net,
    a_x_b_8 => mult7_p_net,
    a_x_b_9 => mult8_p_net,
    a_x_b_10 => mult9_p_net,
    a_x_b_11 => mult10_p_net,
    a_x_b_12 => mult11_p_net,
    a_x_b_13 => mult12_p_net,
    a_x_b_14 => mult13_p_net,
    a_x_b_15 => mult14_p_net,
    a_x_b_16 => mult15_p_net
  );
  vector_reinterpret1 : entity xil_defaultlib.psb3_0_vector_reinterpret1 
  port map (
    in_1 => slice0_y_net_x4,
    in_2 => slice1_y_net_x4,
    in_3 => slice2_y_net_x4,
    in_4 => slice3_y_net_x4,
    in_5 => slice4_y_net_x4,
    in_6 => slice5_y_net_x4,
    in_7 => slice6_y_net_x4,
    in_8 => slice7_y_net_x4,
    in_9 => slice8_y_net_x4,
    in_10 => slice9_y_net_x4,
    in_11 => slice10_y_net_x4,
    in_12 => slice11_y_net_x4,
    in_13 => slice12_y_net_x4,
    in_14 => slice13_y_net_x4,
    in_15 => slice14_y_net_x4,
    in_16 => slice15_y_net_x4,
    out_1 => reinterpret0_output_port_net_x13,
    out_2 => reinterpret1_output_port_net_x13,
    out_3 => reinterpret2_output_port_net_x13,
    out_4 => reinterpret3_output_port_net_x13,
    out_5 => reinterpret4_output_port_net_x13,
    out_6 => reinterpret5_output_port_net_x13,
    out_7 => reinterpret6_output_port_net_x13,
    out_8 => reinterpret7_output_port_net_x13,
    out_9 => reinterpret8_output_port_net_x13,
    out_10 => reinterpret9_output_port_net_x13,
    out_11 => reinterpret10_output_port_net_x13,
    out_12 => reinterpret11_output_port_net_x13,
    out_13 => reinterpret12_output_port_net_x13,
    out_14 => reinterpret13_output_port_net_x13,
    out_15 => reinterpret14_output_port_net_x13,
    out_16 => reinterpret15_output_port_net_x13
  );
  vector_reinterpret10 : entity xil_defaultlib.psb3_0_vector_reinterpret10 
  port map (
    in_1 => slice0_y_net_x2,
    in_2 => slice1_y_net_x2,
    in_3 => slice2_y_net_x2,
    in_4 => slice3_y_net_x2,
    in_5 => slice4_y_net_x2,
    in_6 => slice5_y_net_x2,
    in_7 => slice6_y_net_x2,
    in_8 => slice7_y_net_x2,
    in_9 => slice8_y_net_x2,
    in_10 => slice9_y_net_x2,
    in_11 => slice10_y_net_x2,
    in_12 => slice11_y_net_x2,
    in_13 => slice12_y_net_x2,
    in_14 => slice13_y_net_x2,
    in_15 => slice14_y_net_x2,
    in_16 => slice15_y_net_x2,
    out_1 => reinterpret0_output_port_net_x12,
    out_2 => reinterpret1_output_port_net_x12,
    out_3 => reinterpret2_output_port_net_x12,
    out_4 => reinterpret3_output_port_net_x12,
    out_5 => reinterpret4_output_port_net_x12,
    out_6 => reinterpret5_output_port_net_x12,
    out_7 => reinterpret6_output_port_net_x12,
    out_8 => reinterpret7_output_port_net_x12,
    out_9 => reinterpret8_output_port_net_x12,
    out_10 => reinterpret9_output_port_net_x12,
    out_11 => reinterpret10_output_port_net_x12,
    out_12 => reinterpret11_output_port_net_x12,
    out_13 => reinterpret12_output_port_net_x12,
    out_14 => reinterpret13_output_port_net_x12,
    out_15 => reinterpret14_output_port_net_x12,
    out_16 => reinterpret15_output_port_net_x12
  );
  vector_reinterpret11 : entity xil_defaultlib.psb3_0_vector_reinterpret11 
  port map (
    in_1 => slice0_y_net_x1,
    in_2 => slice1_y_net_x1,
    in_3 => slice2_y_net_x1,
    in_4 => slice3_y_net_x1,
    in_5 => slice4_y_net_x1,
    in_6 => slice5_y_net_x1,
    in_7 => slice6_y_net_x1,
    in_8 => slice7_y_net_x1,
    in_9 => slice8_y_net_x1,
    in_10 => slice9_y_net_x1,
    in_11 => slice10_y_net_x1,
    in_12 => slice11_y_net_x1,
    in_13 => slice12_y_net_x1,
    in_14 => slice13_y_net_x1,
    in_15 => slice14_y_net_x1,
    in_16 => slice15_y_net_x1,
    out_1 => reinterpret0_output_port_net_x11,
    out_2 => reinterpret1_output_port_net_x11,
    out_3 => reinterpret2_output_port_net_x11,
    out_4 => reinterpret3_output_port_net_x11,
    out_5 => reinterpret4_output_port_net_x11,
    out_6 => reinterpret5_output_port_net_x11,
    out_7 => reinterpret6_output_port_net_x11,
    out_8 => reinterpret7_output_port_net_x11,
    out_9 => reinterpret8_output_port_net_x11,
    out_10 => reinterpret9_output_port_net_x11,
    out_11 => reinterpret10_output_port_net_x11,
    out_12 => reinterpret11_output_port_net_x11,
    out_13 => reinterpret12_output_port_net_x11,
    out_14 => reinterpret13_output_port_net_x11,
    out_15 => reinterpret14_output_port_net_x11,
    out_16 => reinterpret15_output_port_net_x11
  );
  vector_reinterpret12 : entity xil_defaultlib.psb3_0_vector_reinterpret12 
  port map (
    in_1 => addsub0_s_net_x2,
    in_2 => addsub1_s_net_x2,
    in_3 => addsub2_s_net_x2,
    in_4 => addsub3_s_net_x2,
    in_5 => addsub4_s_net_x2,
    in_6 => addsub5_s_net_x2,
    in_7 => addsub6_s_net_x1,
    in_8 => addsub7_s_net_x2,
    in_9 => addsub8_s_net_x2,
    in_10 => addsub9_s_net_x2,
    in_11 => addsub10_s_net_x2,
    in_12 => addsub11_s_net_x2,
    in_13 => addsub12_s_net_x2,
    in_14 => addsub13_s_net_x2,
    in_15 => addsub14_s_net_x2,
    in_16 => addsub15_s_net_x2,
    out_1 => reinterpret0_output_port_net_x10,
    out_2 => reinterpret1_output_port_net_x10,
    out_3 => reinterpret2_output_port_net_x10,
    out_4 => reinterpret3_output_port_net_x10,
    out_5 => reinterpret4_output_port_net_x10,
    out_6 => reinterpret5_output_port_net_x10,
    out_7 => reinterpret6_output_port_net_x10,
    out_8 => reinterpret7_output_port_net_x10,
    out_9 => reinterpret8_output_port_net_x10,
    out_10 => reinterpret9_output_port_net_x10,
    out_11 => reinterpret10_output_port_net_x10,
    out_12 => reinterpret11_output_port_net_x10,
    out_13 => reinterpret12_output_port_net_x10,
    out_14 => reinterpret13_output_port_net_x10,
    out_15 => reinterpret14_output_port_net_x10,
    out_16 => reinterpret15_output_port_net_x10
  );
  vector_reinterpret13 : entity xil_defaultlib.psb3_0_vector_reinterpret13 
  port map (
    in_1 => addsub0_s_net_x1,
    in_2 => addsub1_s_net_x1,
    in_3 => addsub2_s_net_x1,
    in_4 => addsub3_s_net_x1,
    in_5 => addsub4_s_net_x1,
    in_6 => addsub5_s_net_x1,
    in_7 => addsub6_s_net_x6,
    in_8 => addsub7_s_net_x1,
    in_9 => addsub8_s_net_x1,
    in_10 => addsub9_s_net_x1,
    in_11 => addsub10_s_net_x1,
    in_12 => addsub11_s_net_x1,
    in_13 => addsub12_s_net_x1,
    in_14 => addsub13_s_net_x1,
    in_15 => addsub14_s_net_x1,
    in_16 => addsub15_s_net_x1,
    out_1 => reinterpret0_output_port_net_x9,
    out_2 => reinterpret1_output_port_net_x9,
    out_3 => reinterpret2_output_port_net_x9,
    out_4 => reinterpret3_output_port_net_x9,
    out_5 => reinterpret4_output_port_net_x9,
    out_6 => reinterpret5_output_port_net_x9,
    out_7 => reinterpret6_output_port_net_x9,
    out_8 => reinterpret7_output_port_net_x9,
    out_9 => reinterpret8_output_port_net_x9,
    out_10 => reinterpret9_output_port_net_x9,
    out_11 => reinterpret10_output_port_net_x9,
    out_12 => reinterpret11_output_port_net_x9,
    out_13 => reinterpret12_output_port_net_x9,
    out_14 => reinterpret13_output_port_net_x9,
    out_15 => reinterpret14_output_port_net_x9,
    out_16 => reinterpret15_output_port_net_x9
  );
  vector_reinterpret14 : entity xil_defaultlib.psb3_0_vector_reinterpret14 
  port map (
    in_1 => slice0_y_net,
    in_2 => slice1_y_net,
    in_3 => slice2_y_net,
    in_4 => slice3_y_net,
    in_5 => slice4_y_net,
    in_6 => slice5_y_net,
    in_7 => slice6_y_net,
    in_8 => slice7_y_net,
    in_9 => slice8_y_net,
    in_10 => slice9_y_net,
    in_11 => slice10_y_net,
    in_12 => slice11_y_net,
    in_13 => slice12_y_net,
    in_14 => slice13_y_net,
    in_15 => slice14_y_net,
    in_16 => slice15_y_net,
    out_1 => reinterpret0_output_port_net_x8,
    out_2 => reinterpret1_output_port_net_x8,
    out_3 => reinterpret2_output_port_net_x8,
    out_4 => reinterpret3_output_port_net_x8,
    out_5 => reinterpret4_output_port_net_x8,
    out_6 => reinterpret5_output_port_net_x8,
    out_7 => reinterpret6_output_port_net_x8,
    out_8 => reinterpret7_output_port_net_x8,
    out_9 => reinterpret8_output_port_net_x8,
    out_10 => reinterpret9_output_port_net_x8,
    out_11 => reinterpret10_output_port_net_x8,
    out_12 => reinterpret11_output_port_net_x8,
    out_13 => reinterpret12_output_port_net_x8,
    out_14 => reinterpret13_output_port_net_x8,
    out_15 => reinterpret14_output_port_net_x8,
    out_16 => reinterpret15_output_port_net_x8
  );
  vector_reinterpret15 : entity xil_defaultlib.psb3_0_vector_reinterpret15 
  port map (
    in_1 => addsub0_s_net_x0,
    in_2 => addsub1_s_net_x0,
    in_3 => addsub2_s_net_x0,
    in_4 => addsub3_s_net_x0,
    in_5 => addsub4_s_net_x0,
    in_6 => addsub5_s_net_x0,
    in_7 => addsub6_s_net_x0,
    in_8 => addsub7_s_net_x0,
    in_9 => addsub8_s_net_x0,
    in_10 => addsub9_s_net_x0,
    in_11 => addsub10_s_net_x0,
    in_12 => addsub11_s_net_x0,
    in_13 => addsub12_s_net_x0,
    in_14 => addsub13_s_net_x0,
    in_15 => addsub14_s_net_x0,
    in_16 => addsub15_s_net_x0,
    out_1 => reinterpret0_output_port_net_x7,
    out_2 => reinterpret1_output_port_net_x7,
    out_3 => reinterpret2_output_port_net_x7,
    out_4 => reinterpret3_output_port_net_x7,
    out_5 => reinterpret4_output_port_net_x7,
    out_6 => reinterpret5_output_port_net_x7,
    out_7 => reinterpret6_output_port_net_x7,
    out_8 => reinterpret7_output_port_net_x7,
    out_9 => reinterpret8_output_port_net_x7,
    out_10 => reinterpret9_output_port_net_x7,
    out_11 => reinterpret10_output_port_net_x7,
    out_12 => reinterpret11_output_port_net_x7,
    out_13 => reinterpret12_output_port_net_x7,
    out_14 => reinterpret13_output_port_net_x7,
    out_15 => reinterpret14_output_port_net_x7,
    out_16 => reinterpret15_output_port_net_x7
  );
  vector_reinterpret16 : entity xil_defaultlib.psb3_0_vector_reinterpret16 
  port map (
    in_1 => addsub0_s_net,
    in_2 => addsub1_s_net,
    in_3 => addsub2_s_net,
    in_4 => addsub3_s_net,
    in_5 => addsub4_s_net,
    in_6 => addsub5_s_net,
    in_7 => addsub6_s_net,
    in_8 => addsub7_s_net,
    in_9 => addsub8_s_net,
    in_10 => addsub9_s_net,
    in_11 => addsub10_s_net,
    in_12 => addsub11_s_net,
    in_13 => addsub12_s_net,
    in_14 => addsub13_s_net,
    in_15 => addsub14_s_net,
    in_16 => addsub15_s_net,
    out_1 => reinterpret0_output_port_net_x6,
    out_2 => reinterpret1_output_port_net_x6,
    out_3 => reinterpret2_output_port_net_x6,
    out_4 => reinterpret3_output_port_net_x6,
    out_5 => reinterpret4_output_port_net_x6,
    out_6 => reinterpret5_output_port_net_x6,
    out_7 => reinterpret6_output_port_net_x6,
    out_8 => reinterpret7_output_port_net_x6,
    out_9 => reinterpret8_output_port_net_x6,
    out_10 => reinterpret9_output_port_net_x6,
    out_11 => reinterpret10_output_port_net_x6,
    out_12 => reinterpret11_output_port_net_x6,
    out_13 => reinterpret12_output_port_net_x6,
    out_14 => reinterpret13_output_port_net_x6,
    out_15 => reinterpret14_output_port_net_x6,
    out_16 => reinterpret15_output_port_net_x6
  );
  vector_reinterpret2 : entity xil_defaultlib.psb3_0_vector_reinterpret2 
  port map (
    in_1 => slice0_y_net_x6,
    in_2 => slice1_y_net_x6,
    in_3 => slice2_y_net_x6,
    in_4 => slice3_y_net_x6,
    in_5 => slice4_y_net_x6,
    in_6 => slice5_y_net_x6,
    in_7 => slice6_y_net_x6,
    in_8 => slice7_y_net_x6,
    in_9 => slice8_y_net_x6,
    in_10 => slice9_y_net_x6,
    in_11 => slice10_y_net_x6,
    in_12 => slice11_y_net_x6,
    in_13 => slice12_y_net_x6,
    in_14 => slice13_y_net_x6,
    in_15 => slice14_y_net_x6,
    in_16 => slice15_y_net_x6,
    out_1 => reinterpret0_output_port_net_x5,
    out_2 => reinterpret1_output_port_net_x5,
    out_3 => reinterpret2_output_port_net_x5,
    out_4 => reinterpret3_output_port_net_x5,
    out_5 => reinterpret4_output_port_net_x5,
    out_6 => reinterpret5_output_port_net_x5,
    out_7 => reinterpret6_output_port_net_x5,
    out_8 => reinterpret7_output_port_net_x5,
    out_9 => reinterpret8_output_port_net_x5,
    out_10 => reinterpret9_output_port_net_x5,
    out_11 => reinterpret10_output_port_net_x5,
    out_12 => reinterpret11_output_port_net_x5,
    out_13 => reinterpret12_output_port_net_x5,
    out_14 => reinterpret13_output_port_net_x5,
    out_15 => reinterpret14_output_port_net_x5,
    out_16 => reinterpret15_output_port_net_x5
  );
  vector_reinterpret3 : entity xil_defaultlib.psb3_0_vector_reinterpret3 
  port map (
    in_1 => slice0_y_net_x5,
    in_2 => slice1_y_net_x5,
    in_3 => slice2_y_net_x5,
    in_4 => slice3_y_net_x5,
    in_5 => slice4_y_net_x5,
    in_6 => slice5_y_net_x5,
    in_7 => slice6_y_net_x5,
    in_8 => slice7_y_net_x5,
    in_9 => slice8_y_net_x5,
    in_10 => slice9_y_net_x5,
    in_11 => slice10_y_net_x5,
    in_12 => slice11_y_net_x5,
    in_13 => slice12_y_net_x5,
    in_14 => slice13_y_net_x5,
    in_15 => slice14_y_net_x5,
    in_16 => slice15_y_net_x5,
    out_1 => reinterpret0_output_port_net_x4,
    out_2 => reinterpret1_output_port_net_x4,
    out_3 => reinterpret2_output_port_net_x4,
    out_4 => reinterpret3_output_port_net_x4,
    out_5 => reinterpret4_output_port_net_x4,
    out_6 => reinterpret5_output_port_net_x4,
    out_7 => reinterpret6_output_port_net_x4,
    out_8 => reinterpret7_output_port_net_x4,
    out_9 => reinterpret8_output_port_net_x4,
    out_10 => reinterpret9_output_port_net_x4,
    out_11 => reinterpret10_output_port_net_x4,
    out_12 => reinterpret11_output_port_net_x4,
    out_13 => reinterpret12_output_port_net_x4,
    out_14 => reinterpret13_output_port_net_x4,
    out_15 => reinterpret14_output_port_net_x4,
    out_16 => reinterpret15_output_port_net_x4
  );
  vector_reinterpret4 : entity xil_defaultlib.psb3_0_vector_reinterpret4 
  port map (
    in_1 => addsub0_s_net_x6,
    in_2 => addsub1_s_net_x6,
    in_3 => addsub2_s_net_x6,
    in_4 => addsub3_s_net_x6,
    in_5 => addsub4_s_net_x6,
    in_6 => addsub5_s_net_x6,
    in_7 => addsub6_s_net_x5,
    in_8 => addsub7_s_net_x6,
    in_9 => addsub8_s_net_x6,
    in_10 => addsub9_s_net_x6,
    in_11 => addsub10_s_net_x6,
    in_12 => addsub11_s_net_x6,
    in_13 => addsub12_s_net_x6,
    in_14 => addsub13_s_net_x6,
    in_15 => addsub14_s_net_x6,
    in_16 => addsub15_s_net_x6,
    out_1 => reinterpret0_output_port_net_x3,
    out_2 => reinterpret1_output_port_net_x3,
    out_3 => reinterpret2_output_port_net_x3,
    out_4 => reinterpret3_output_port_net_x3,
    out_5 => reinterpret4_output_port_net_x3,
    out_6 => reinterpret5_output_port_net_x3,
    out_7 => reinterpret6_output_port_net_x3,
    out_8 => reinterpret7_output_port_net_x3,
    out_9 => reinterpret8_output_port_net_x3,
    out_10 => reinterpret9_output_port_net_x3,
    out_11 => reinterpret10_output_port_net_x3,
    out_12 => reinterpret11_output_port_net_x3,
    out_13 => reinterpret12_output_port_net_x3,
    out_14 => reinterpret13_output_port_net_x3,
    out_15 => reinterpret14_output_port_net_x3,
    out_16 => reinterpret15_output_port_net_x3
  );
  vector_reinterpret5 : entity xil_defaultlib.psb3_0_vector_reinterpret5 
  port map (
    in_1 => addsub0_s_net_x5,
    in_2 => addsub1_s_net_x5,
    in_3 => addsub2_s_net_x5,
    in_4 => addsub3_s_net_x5,
    in_5 => addsub4_s_net_x5,
    in_6 => addsub5_s_net_x5,
    in_7 => addsub6_s_net_x4,
    in_8 => addsub7_s_net_x5,
    in_9 => addsub8_s_net_x5,
    in_10 => addsub9_s_net_x5,
    in_11 => addsub10_s_net_x5,
    in_12 => addsub11_s_net_x5,
    in_13 => addsub12_s_net_x5,
    in_14 => addsub13_s_net_x5,
    in_15 => addsub14_s_net_x5,
    in_16 => addsub15_s_net_x5,
    out_1 => reinterpret0_output_port_net_x2,
    out_2 => reinterpret1_output_port_net_x2,
    out_3 => reinterpret2_output_port_net_x2,
    out_4 => reinterpret3_output_port_net_x2,
    out_5 => reinterpret4_output_port_net_x2,
    out_6 => reinterpret5_output_port_net_x2,
    out_7 => reinterpret6_output_port_net_x2,
    out_8 => reinterpret7_output_port_net_x2,
    out_9 => reinterpret8_output_port_net_x2,
    out_10 => reinterpret9_output_port_net_x2,
    out_11 => reinterpret10_output_port_net_x2,
    out_12 => reinterpret11_output_port_net_x2,
    out_13 => reinterpret12_output_port_net_x2,
    out_14 => reinterpret13_output_port_net_x2,
    out_15 => reinterpret14_output_port_net_x2,
    out_16 => reinterpret15_output_port_net_x2
  );
  vector_reinterpret6 : entity xil_defaultlib.psb3_0_vector_reinterpret6 
  port map (
    in_1 => slice0_y_net_x3,
    in_2 => slice1_y_net_x3,
    in_3 => slice2_y_net_x3,
    in_4 => slice3_y_net_x3,
    in_5 => slice4_y_net_x3,
    in_6 => slice5_y_net_x3,
    in_7 => slice6_y_net_x3,
    in_8 => slice7_y_net_x3,
    in_9 => slice8_y_net_x3,
    in_10 => slice9_y_net_x3,
    in_11 => slice10_y_net_x3,
    in_12 => slice11_y_net_x3,
    in_13 => slice12_y_net_x3,
    in_14 => slice13_y_net_x3,
    in_15 => slice14_y_net_x3,
    in_16 => slice15_y_net_x3,
    out_1 => reinterpret0_output_port_net_x1,
    out_2 => reinterpret1_output_port_net_x1,
    out_3 => reinterpret2_output_port_net_x1,
    out_4 => reinterpret3_output_port_net_x1,
    out_5 => reinterpret4_output_port_net_x1,
    out_6 => reinterpret5_output_port_net_x1,
    out_7 => reinterpret6_output_port_net_x1,
    out_8 => reinterpret7_output_port_net_x1,
    out_9 => reinterpret8_output_port_net_x1,
    out_10 => reinterpret9_output_port_net_x1,
    out_11 => reinterpret10_output_port_net_x1,
    out_12 => reinterpret11_output_port_net_x1,
    out_13 => reinterpret12_output_port_net_x1,
    out_14 => reinterpret13_output_port_net_x1,
    out_15 => reinterpret14_output_port_net_x1,
    out_16 => reinterpret15_output_port_net_x1
  );
  vector_reinterpret7 : entity xil_defaultlib.psb3_0_vector_reinterpret7 
  port map (
    in_1 => addsub0_s_net_x4,
    in_2 => addsub1_s_net_x4,
    in_3 => addsub2_s_net_x4,
    in_4 => addsub3_s_net_x4,
    in_5 => addsub4_s_net_x4,
    in_6 => addsub5_s_net_x4,
    in_7 => addsub6_s_net_x3,
    in_8 => addsub7_s_net_x4,
    in_9 => addsub8_s_net_x4,
    in_10 => addsub9_s_net_x4,
    in_11 => addsub10_s_net_x4,
    in_12 => addsub11_s_net_x4,
    in_13 => addsub12_s_net_x4,
    in_14 => addsub13_s_net_x4,
    in_15 => addsub14_s_net_x4,
    in_16 => addsub15_s_net_x4,
    out_1 => reinterpret0_output_port_net_x0,
    out_2 => reinterpret1_output_port_net_x0,
    out_3 => reinterpret2_output_port_net_x0,
    out_4 => reinterpret3_output_port_net_x0,
    out_5 => reinterpret4_output_port_net_x0,
    out_6 => reinterpret5_output_port_net_x0,
    out_7 => reinterpret6_output_port_net_x0,
    out_8 => reinterpret7_output_port_net_x0,
    out_9 => reinterpret8_output_port_net_x0,
    out_10 => reinterpret9_output_port_net_x0,
    out_11 => reinterpret10_output_port_net_x0,
    out_12 => reinterpret11_output_port_net_x0,
    out_13 => reinterpret12_output_port_net_x0,
    out_14 => reinterpret13_output_port_net_x0,
    out_15 => reinterpret14_output_port_net_x0,
    out_16 => reinterpret15_output_port_net_x0
  );
  vector_reinterpret8 : entity xil_defaultlib.psb3_0_vector_reinterpret8 
  port map (
    in_1 => addsub0_s_net_x3,
    in_2 => addsub1_s_net_x3,
    in_3 => addsub2_s_net_x3,
    in_4 => addsub3_s_net_x3,
    in_5 => addsub4_s_net_x3,
    in_6 => addsub5_s_net_x3,
    in_7 => addsub6_s_net_x2,
    in_8 => addsub7_s_net_x3,
    in_9 => addsub8_s_net_x3,
    in_10 => addsub9_s_net_x3,
    in_11 => addsub10_s_net_x3,
    in_12 => addsub11_s_net_x3,
    in_13 => addsub12_s_net_x3,
    in_14 => addsub13_s_net_x3,
    in_15 => addsub14_s_net_x3,
    in_16 => addsub15_s_net_x3,
    out_1 => reinterpret0_output_port_net,
    out_2 => reinterpret1_output_port_net,
    out_3 => reinterpret2_output_port_net,
    out_4 => reinterpret3_output_port_net,
    out_5 => reinterpret4_output_port_net,
    out_6 => reinterpret5_output_port_net,
    out_7 => reinterpret6_output_port_net,
    out_8 => reinterpret7_output_port_net,
    out_9 => reinterpret8_output_port_net,
    out_10 => reinterpret9_output_port_net,
    out_11 => reinterpret10_output_port_net,
    out_12 => reinterpret11_output_port_net,
    out_13 => reinterpret12_output_port_net,
    out_14 => reinterpret13_output_port_net,
    out_15 => reinterpret14_output_port_net,
    out_16 => reinterpret15_output_port_net
  );
  vector_reinterpret9 : entity xil_defaultlib.psb3_0_vector_reinterpret9 
  port map (
    in_1 => slice0_y_net_x0,
    in_2 => slice1_y_net_x0,
    in_3 => slice2_y_net_x0,
    in_4 => slice3_y_net_x0,
    in_5 => slice4_y_net_x0,
    in_6 => slice5_y_net_x0,
    in_7 => slice6_y_net_x0,
    in_8 => slice7_y_net_x0,
    in_9 => slice8_y_net_x0,
    in_10 => slice9_y_net_x0,
    in_11 => slice10_y_net_x0,
    in_12 => slice11_y_net_x0,
    in_13 => slice12_y_net_x0,
    in_14 => slice13_y_net_x0,
    in_15 => slice14_y_net_x0,
    in_16 => slice15_y_net_x0,
    out_1 => reinterpret0_output_port_net_x26,
    out_2 => reinterpret1_output_port_net_x27,
    out_3 => reinterpret2_output_port_net_x27,
    out_4 => reinterpret3_output_port_net_x27,
    out_5 => reinterpret4_output_port_net_x27,
    out_6 => reinterpret5_output_port_net_x27,
    out_7 => reinterpret6_output_port_net_x27,
    out_8 => reinterpret7_output_port_net_x27,
    out_9 => reinterpret8_output_port_net_x26,
    out_10 => reinterpret9_output_port_net_x26,
    out_11 => reinterpret10_output_port_net_x26,
    out_12 => reinterpret11_output_port_net_x26,
    out_13 => reinterpret12_output_port_net_x26,
    out_14 => reinterpret13_output_port_net_x26,
    out_15 => reinterpret14_output_port_net_x26,
    out_16 => reinterpret15_output_port_net_x26
  );
  vector_to_scalar : entity xil_defaultlib.psb3_0_vector_to_scalar_x7 
  port map (
    i_1 => reinterpret0_output_port_net_x3,
    i_2 => reinterpret1_output_port_net_x3,
    i_3 => reinterpret2_output_port_net_x3,
    i_4 => reinterpret3_output_port_net_x3,
    i_5 => reinterpret4_output_port_net_x3,
    i_6 => reinterpret5_output_port_net_x3,
    i_7 => reinterpret6_output_port_net_x3,
    i_8 => reinterpret7_output_port_net_x3,
    i_9 => reinterpret8_output_port_net_x3,
    i_10 => reinterpret9_output_port_net_x3,
    i_11 => reinterpret10_output_port_net_x3,
    i_12 => reinterpret11_output_port_net_x3,
    i_13 => reinterpret12_output_port_net_x3,
    i_14 => reinterpret13_output_port_net_x3,
    i_15 => reinterpret14_output_port_net_x3,
    i_16 => reinterpret15_output_port_net_x3,
    o => concat1_y_net_x6
  );
  vector_to_scalar1 : entity xil_defaultlib.psb3_0_vector_to_scalar1_x7 
  port map (
    i_1 => reinterpret0_output_port_net_x2,
    i_2 => reinterpret1_output_port_net_x2,
    i_3 => reinterpret2_output_port_net_x2,
    i_4 => reinterpret3_output_port_net_x2,
    i_5 => reinterpret4_output_port_net_x2,
    i_6 => reinterpret5_output_port_net_x2,
    i_7 => reinterpret6_output_port_net_x2,
    i_8 => reinterpret7_output_port_net_x2,
    i_9 => reinterpret8_output_port_net_x2,
    i_10 => reinterpret9_output_port_net_x2,
    i_11 => reinterpret10_output_port_net_x2,
    i_12 => reinterpret11_output_port_net_x2,
    i_13 => reinterpret12_output_port_net_x2,
    i_14 => reinterpret13_output_port_net_x2,
    i_15 => reinterpret14_output_port_net_x2,
    i_16 => reinterpret15_output_port_net_x2,
    o => concat1_y_net_x5
  );
  vector_to_scalar2 : entity xil_defaultlib.psb3_0_vector_to_scalar2_x7 
  port map (
    i_1 => reinterpret0_output_port_net_x0,
    i_2 => reinterpret1_output_port_net_x0,
    i_3 => reinterpret2_output_port_net_x0,
    i_4 => reinterpret3_output_port_net_x0,
    i_5 => reinterpret4_output_port_net_x0,
    i_6 => reinterpret5_output_port_net_x0,
    i_7 => reinterpret6_output_port_net_x0,
    i_8 => reinterpret7_output_port_net_x0,
    i_9 => reinterpret8_output_port_net_x0,
    i_10 => reinterpret9_output_port_net_x0,
    i_11 => reinterpret10_output_port_net_x0,
    i_12 => reinterpret11_output_port_net_x0,
    i_13 => reinterpret12_output_port_net_x0,
    i_14 => reinterpret13_output_port_net_x0,
    i_15 => reinterpret14_output_port_net_x0,
    i_16 => reinterpret15_output_port_net_x0,
    o => concat1_y_net_x4
  );
  vector_to_scalar3 : entity xil_defaultlib.psb3_0_vector_to_scalar3 
  port map (
    i_1 => reinterpret0_output_port_net,
    i_2 => reinterpret1_output_port_net,
    i_3 => reinterpret2_output_port_net,
    i_4 => reinterpret3_output_port_net,
    i_5 => reinterpret4_output_port_net,
    i_6 => reinterpret5_output_port_net,
    i_7 => reinterpret6_output_port_net,
    i_8 => reinterpret7_output_port_net,
    i_9 => reinterpret8_output_port_net,
    i_10 => reinterpret9_output_port_net,
    i_11 => reinterpret10_output_port_net,
    i_12 => reinterpret11_output_port_net,
    i_13 => reinterpret12_output_port_net,
    i_14 => reinterpret13_output_port_net,
    i_15 => reinterpret14_output_port_net,
    i_16 => reinterpret15_output_port_net,
    o => concat1_y_net_x3
  );
  vector_to_scalar4 : entity xil_defaultlib.psb3_0_vector_to_scalar4 
  port map (
    i_1 => reinterpret0_output_port_net_x10,
    i_2 => reinterpret1_output_port_net_x10,
    i_3 => reinterpret2_output_port_net_x10,
    i_4 => reinterpret3_output_port_net_x10,
    i_5 => reinterpret4_output_port_net_x10,
    i_6 => reinterpret5_output_port_net_x10,
    i_7 => reinterpret6_output_port_net_x10,
    i_8 => reinterpret7_output_port_net_x10,
    i_9 => reinterpret8_output_port_net_x10,
    i_10 => reinterpret9_output_port_net_x10,
    i_11 => reinterpret10_output_port_net_x10,
    i_12 => reinterpret11_output_port_net_x10,
    i_13 => reinterpret12_output_port_net_x10,
    i_14 => reinterpret13_output_port_net_x10,
    i_15 => reinterpret14_output_port_net_x10,
    i_16 => reinterpret15_output_port_net_x10,
    o => concat1_y_net_x2
  );
  vector_to_scalar5 : entity xil_defaultlib.psb3_0_vector_to_scalar5 
  port map (
    i_1 => reinterpret0_output_port_net_x9,
    i_2 => reinterpret1_output_port_net_x9,
    i_3 => reinterpret2_output_port_net_x9,
    i_4 => reinterpret3_output_port_net_x9,
    i_5 => reinterpret4_output_port_net_x9,
    i_6 => reinterpret5_output_port_net_x9,
    i_7 => reinterpret6_output_port_net_x9,
    i_8 => reinterpret7_output_port_net_x9,
    i_9 => reinterpret8_output_port_net_x9,
    i_10 => reinterpret9_output_port_net_x9,
    i_11 => reinterpret10_output_port_net_x9,
    i_12 => reinterpret11_output_port_net_x9,
    i_13 => reinterpret12_output_port_net_x9,
    i_14 => reinterpret13_output_port_net_x9,
    i_15 => reinterpret14_output_port_net_x9,
    i_16 => reinterpret15_output_port_net_x9,
    o => concat1_y_net_x1
  );
  vector_to_scalar6 : entity xil_defaultlib.psb3_0_vector_to_scalar6 
  port map (
    i_1 => reinterpret0_output_port_net_x7,
    i_2 => reinterpret1_output_port_net_x7,
    i_3 => reinterpret2_output_port_net_x7,
    i_4 => reinterpret3_output_port_net_x7,
    i_5 => reinterpret4_output_port_net_x7,
    i_6 => reinterpret5_output_port_net_x7,
    i_7 => reinterpret6_output_port_net_x7,
    i_8 => reinterpret7_output_port_net_x7,
    i_9 => reinterpret8_output_port_net_x7,
    i_10 => reinterpret9_output_port_net_x7,
    i_11 => reinterpret10_output_port_net_x7,
    i_12 => reinterpret11_output_port_net_x7,
    i_13 => reinterpret12_output_port_net_x7,
    i_14 => reinterpret13_output_port_net_x7,
    i_15 => reinterpret14_output_port_net_x7,
    i_16 => reinterpret15_output_port_net_x7,
    o => concat1_y_net_x0
  );
  vector_to_scalar7 : entity xil_defaultlib.psb3_0_vector_to_scalar7 
  port map (
    i_1 => reinterpret0_output_port_net_x6,
    i_2 => reinterpret1_output_port_net_x6,
    i_3 => reinterpret2_output_port_net_x6,
    i_4 => reinterpret3_output_port_net_x6,
    i_5 => reinterpret4_output_port_net_x6,
    i_6 => reinterpret5_output_port_net_x6,
    i_7 => reinterpret6_output_port_net_x6,
    i_8 => reinterpret7_output_port_net_x6,
    i_9 => reinterpret8_output_port_net_x6,
    i_10 => reinterpret9_output_port_net_x6,
    i_11 => reinterpret10_output_port_net_x6,
    i_12 => reinterpret11_output_port_net_x6,
    i_13 => reinterpret12_output_port_net_x6,
    i_14 => reinterpret13_output_port_net_x6,
    i_15 => reinterpret14_output_port_net_x6,
    i_16 => reinterpret15_output_port_net_x6,
    o => concat1_y_net
  );
  delaycounter : entity xil_defaultlib.psb3_0_delaycounter 
  port map (
    edge1 => delay11_q_net,
    edge2 => test_systolicfft_vhdl_black_box_vo_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    delay => counter1_op_net_x7
  );
  ov_detector_ifft_im : entity xil_defaultlib.psb3_0_ov_detector_ifft_im 
  port map (
    rst => gin_tl_reset_net,
    a_1 => reinterpret16_output_port_net,
    b_1 => mux0_y_net,
    en => test_systolicfft_vhdl_black_box_vo_net,
    a_2 => reinterpret17_output_port_net,
    a_3 => reinterpret18_output_port_net,
    a_4 => reinterpret19_output_port_net,
    a_5 => reinterpret20_output_port_net,
    a_6 => reinterpret21_output_port_net,
    a_7 => reinterpret22_output_port_net,
    a_8 => reinterpret23_output_port_net,
    b_2 => mux1_y_net,
    b_3 => mux2_y_net,
    b_4 => mux3_y_net,
    b_5 => mux4_y_net,
    b_6 => mux5_y_net,
    b_7 => mux6_y_net,
    b_8 => mux7_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    ov => register_q_net_x9
  );
  ov_detector_ifft_re : entity xil_defaultlib.psb3_0_ov_detector_ifft_re 
  port map (
    rst => gin_tl_reset_net,
    a_1 => reinterpret24_output_port_net,
    b_1 => mux0_y_net_x0,
    en => test_systolicfft_vhdl_black_box_vo_net,
    a_2 => reinterpret25_output_port_net,
    a_3 => reinterpret26_output_port_net,
    a_4 => reinterpret27_output_port_net,
    a_5 => reinterpret28_output_port_net,
    a_6 => reinterpret29_output_port_net,
    a_7 => reinterpret30_output_port_net,
    a_8 => reinterpret31_output_port_net,
    b_2 => mux1_y_net_x0,
    b_3 => mux2_y_net_x0,
    b_4 => mux3_y_net_x0,
    b_5 => mux4_y_net_x0,
    b_6 => mux5_y_net_x0,
    b_7 => mux6_y_net_x0,
    b_8 => mux7_y_net_x0,
    clk_1 => clk_net,
    ce_1 => ce_net,
    ov => register_q_net_x8
  );
  reordering_extending_buffer_imag_1 : entity xil_defaultlib.psb3_0_reordering_extending_buffer_imag_1 
  port map (
    in_reset => gin_tl_reset_net,
    input1 => mux0_y_net,
    input2 => mux4_y_net,
    in_tvalid => delay19_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    vec_output_1 => reinterpret0_output_port_net_x25,
    vec_output_2 => reinterpret1_output_port_net_x26,
    vec_output_3 => reinterpret2_output_port_net_x26,
    vec_output_4 => reinterpret3_output_port_net_x26,
    vec_output_5 => reinterpret4_output_port_net_x26,
    vec_output_6 => reinterpret5_output_port_net_x26,
    vec_output_7 => reinterpret6_output_port_net_x26,
    vec_output_8 => reinterpret7_output_port_net_x26,
    vec_output_9 => reinterpret8_output_port_net_x25,
    vec_output_10 => reinterpret9_output_port_net_x25,
    vec_output_11 => reinterpret10_output_port_net_x25,
    vec_output_12 => reinterpret11_output_port_net_x25,
    vec_output_13 => reinterpret12_output_port_net_x25,
    vec_output_14 => reinterpret13_output_port_net_x25,
    vec_output_15 => reinterpret14_output_port_net_x25,
    vec_output_16 => reinterpret15_output_port_net_x25
  );
  reordering_extending_buffer_imag_2 : entity xil_defaultlib.psb3_0_reordering_extending_buffer_imag_2 
  port map (
    in_reset => gin_tl_reset_net,
    input1 => mux1_y_net,
    input2 => mux5_y_net,
    in_tvalid => delay19_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    vec_output_1 => reinterpret0_output_port_net_x24,
    vec_output_2 => reinterpret1_output_port_net_x25,
    vec_output_3 => reinterpret2_output_port_net_x25,
    vec_output_4 => reinterpret3_output_port_net_x25,
    vec_output_5 => reinterpret4_output_port_net_x25,
    vec_output_6 => reinterpret5_output_port_net_x25,
    vec_output_7 => reinterpret6_output_port_net_x25,
    vec_output_8 => reinterpret7_output_port_net_x25,
    vec_output_9 => reinterpret8_output_port_net_x14,
    vec_output_10 => reinterpret9_output_port_net_x24,
    vec_output_11 => reinterpret10_output_port_net_x24,
    vec_output_12 => reinterpret11_output_port_net_x24,
    vec_output_13 => reinterpret12_output_port_net_x24,
    vec_output_14 => reinterpret13_output_port_net_x24,
    vec_output_15 => reinterpret14_output_port_net_x24,
    vec_output_16 => reinterpret15_output_port_net_x24
  );
  reordering_extending_buffer_imag_3 : entity xil_defaultlib.psb3_0_reordering_extending_buffer_imag_3 
  port map (
    in_reset => gin_tl_reset_net,
    input1 => mux2_y_net,
    input2 => mux6_y_net,
    in_tvalid => delay19_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    vec_output_1 => reinterpret0_output_port_net_x23,
    vec_output_2 => reinterpret1_output_port_net_x24,
    vec_output_3 => reinterpret2_output_port_net_x24,
    vec_output_4 => reinterpret3_output_port_net_x24,
    vec_output_5 => reinterpret4_output_port_net_x24,
    vec_output_6 => reinterpret5_output_port_net_x24,
    vec_output_7 => reinterpret6_output_port_net_x24,
    vec_output_8 => reinterpret7_output_port_net_x24,
    vec_output_9 => reinterpret8_output_port_net_x24,
    vec_output_10 => reinterpret9_output_port_net_x23,
    vec_output_11 => reinterpret10_output_port_net_x23,
    vec_output_12 => reinterpret11_output_port_net_x23,
    vec_output_13 => reinterpret12_output_port_net_x23,
    vec_output_14 => reinterpret13_output_port_net_x23,
    vec_output_15 => reinterpret14_output_port_net_x23,
    vec_output_16 => reinterpret15_output_port_net_x23
  );
  reordering_extending_buffer_imag_4 : entity xil_defaultlib.psb3_0_reordering_extending_buffer_imag_4 
  port map (
    in_reset => gin_tl_reset_net,
    input1 => mux3_y_net,
    input2 => mux7_y_net,
    in_tvalid => delay19_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    vec_output_1 => reinterpret0_output_port_net_x22,
    vec_output_2 => reinterpret1_output_port_net_x23,
    vec_output_3 => reinterpret2_output_port_net_x23,
    vec_output_4 => reinterpret3_output_port_net_x23,
    vec_output_5 => reinterpret4_output_port_net_x23,
    vec_output_6 => reinterpret5_output_port_net_x23,
    vec_output_7 => reinterpret6_output_port_net_x23,
    vec_output_8 => reinterpret7_output_port_net_x23,
    vec_output_9 => reinterpret8_output_port_net_x23,
    vec_output_10 => reinterpret9_output_port_net_x22,
    vec_output_11 => reinterpret10_output_port_net_x22,
    vec_output_12 => reinterpret11_output_port_net_x22,
    vec_output_13 => reinterpret12_output_port_net_x22,
    vec_output_14 => reinterpret13_output_port_net_x22,
    vec_output_15 => reinterpret14_output_port_net_x22,
    vec_output_16 => reinterpret15_output_port_net_x22
  );
  reordering_extending_buffer_real_1 : entity xil_defaultlib.psb3_0_reordering_extending_buffer_real_1 
  port map (
    in_reset => gin_tl_reset_net,
    input1 => mux0_y_net_x0,
    input2 => mux4_y_net_x0,
    in_tvalid => delay19_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    vec_output_1 => reinterpret0_output_port_net_x21,
    out_tvalid => delay8_q_net_x3,
    vec_output_2 => reinterpret1_output_port_net_x22,
    vec_output_3 => reinterpret2_output_port_net_x22,
    vec_output_4 => reinterpret3_output_port_net_x22,
    vec_output_5 => reinterpret4_output_port_net_x22,
    vec_output_6 => reinterpret5_output_port_net_x22,
    vec_output_7 => reinterpret6_output_port_net_x22,
    vec_output_8 => reinterpret7_output_port_net_x22,
    vec_output_9 => reinterpret8_output_port_net_x22,
    vec_output_10 => reinterpret9_output_port_net_x21,
    vec_output_11 => reinterpret10_output_port_net_x21,
    vec_output_12 => reinterpret11_output_port_net_x21,
    vec_output_13 => reinterpret12_output_port_net_x21,
    vec_output_14 => reinterpret13_output_port_net_x21,
    vec_output_15 => reinterpret14_output_port_net_x21,
    vec_output_16 => reinterpret15_output_port_net_x21
  );
  reordering_extending_buffer_real_2 : entity xil_defaultlib.psb3_0_reordering_extending_buffer_real_2 
  port map (
    in_reset => gin_tl_reset_net,
    input1 => mux1_y_net_x0,
    input2 => mux5_y_net_x0,
    in_tvalid => delay19_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    vec_output_1 => reinterpret0_output_port_net_x20,
    vec_output_2 => reinterpret1_output_port_net_x21,
    vec_output_3 => reinterpret2_output_port_net_x21,
    vec_output_4 => reinterpret3_output_port_net_x21,
    vec_output_5 => reinterpret4_output_port_net_x21,
    vec_output_6 => reinterpret5_output_port_net_x21,
    vec_output_7 => reinterpret6_output_port_net_x21,
    vec_output_8 => reinterpret7_output_port_net_x21,
    vec_output_9 => reinterpret8_output_port_net_x21,
    vec_output_10 => reinterpret9_output_port_net_x20,
    vec_output_11 => reinterpret10_output_port_net_x20,
    vec_output_12 => reinterpret11_output_port_net_x20,
    vec_output_13 => reinterpret12_output_port_net_x20,
    vec_output_14 => reinterpret13_output_port_net_x20,
    vec_output_15 => reinterpret14_output_port_net_x20,
    vec_output_16 => reinterpret15_output_port_net_x20
  );
  reordering_extending_buffer_real_3 : entity xil_defaultlib.psb3_0_reordering_extending_buffer_real_3 
  port map (
    in_reset => gin_tl_reset_net,
    input1 => mux2_y_net_x0,
    input2 => mux6_y_net_x0,
    in_tvalid => delay19_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    vec_output_1 => reinterpret0_output_port_net_x19,
    vec_output_2 => reinterpret1_output_port_net_x20,
    vec_output_3 => reinterpret2_output_port_net_x20,
    vec_output_4 => reinterpret3_output_port_net_x20,
    vec_output_5 => reinterpret4_output_port_net_x20,
    vec_output_6 => reinterpret5_output_port_net_x20,
    vec_output_7 => reinterpret6_output_port_net_x20,
    vec_output_8 => reinterpret7_output_port_net_x20,
    vec_output_9 => reinterpret8_output_port_net_x20,
    vec_output_10 => reinterpret9_output_port_net_x19,
    vec_output_11 => reinterpret10_output_port_net_x19,
    vec_output_12 => reinterpret11_output_port_net_x19,
    vec_output_13 => reinterpret12_output_port_net_x19,
    vec_output_14 => reinterpret13_output_port_net_x19,
    vec_output_15 => reinterpret14_output_port_net_x19,
    vec_output_16 => reinterpret15_output_port_net_x19
  );
  reordering_extending_buffer_real_4 : entity xil_defaultlib.psb3_0_reordering_extending_buffer_real_4 
  port map (
    in_reset => gin_tl_reset_net,
    input1 => mux3_y_net_x0,
    input2 => mux7_y_net_x0,
    in_tvalid => delay19_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    vec_output_1 => reinterpret0_output_port_net_x18,
    vec_output_2 => reinterpret1_output_port_net_x19,
    vec_output_3 => reinterpret2_output_port_net_x19,
    vec_output_4 => reinterpret3_output_port_net_x19,
    vec_output_5 => reinterpret4_output_port_net_x19,
    vec_output_6 => reinterpret5_output_port_net_x19,
    vec_output_7 => reinterpret6_output_port_net_x19,
    vec_output_8 => reinterpret7_output_port_net_x19,
    vec_output_9 => reinterpret8_output_port_net_x19,
    vec_output_10 => reinterpret9_output_port_net_x18,
    vec_output_11 => reinterpret10_output_port_net_x18,
    vec_output_12 => reinterpret11_output_port_net_x18,
    vec_output_13 => reinterpret12_output_port_net_x18,
    vec_output_14 => reinterpret13_output_port_net_x18,
    vec_output_15 => reinterpret14_output_port_net_x18,
    vec_output_16 => reinterpret15_output_port_net_x18
  );
  vector_ifft : entity xil_defaultlib.psb3_0_vector_ifft 
  port map (
    i_re_1 => mux2_y_net_x1,
    i_im_1 => mux27_y_net,
    vi => delay11_q_net,
    si => constant15_op_net,
    i_re_2 => mux29_y_net,
    i_re_3 => mux33_y_net,
    i_re_4 => mux37_y_net,
    i_re_5 => mux41_y_net,
    i_re_6 => mux45_y_net,
    i_re_7 => mux49_y_net,
    i_re_8 => mux53_y_net,
    i_im_2 => mux30_y_net,
    i_im_3 => mux34_y_net,
    i_im_4 => mux38_y_net,
    i_im_5 => mux42_y_net,
    i_im_6 => mux46_y_net,
    i_im_7 => mux50_y_net,
    i_im_8 => mux54_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    o_re_1 => reinterpret24_output_port_net,
    o_im_1 => reinterpret16_output_port_net,
    vo => test_systolicfft_vhdl_black_box_vo_net,
    o_re_2 => reinterpret25_output_port_net,
    o_re_3 => reinterpret26_output_port_net,
    o_re_4 => reinterpret27_output_port_net,
    o_re_5 => reinterpret28_output_port_net,
    o_re_6 => reinterpret29_output_port_net,
    o_re_7 => reinterpret30_output_port_net,
    o_re_8 => reinterpret31_output_port_net,
    o_im_2 => reinterpret17_output_port_net,
    o_im_3 => reinterpret18_output_port_net,
    o_im_4 => reinterpret19_output_port_net,
    o_im_5 => reinterpret20_output_port_net,
    o_im_6 => reinterpret21_output_port_net,
    o_im_7 => reinterpret22_output_port_net,
    o_im_8 => reinterpret23_output_port_net
  );
  bitbasher1 : entity xil_defaultlib.sysgen_bitbasher_086dfd1ec3 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in_x0 => fifo2_dout_net,
    a => bitbasher1_a_net,
    b => bitbasher1_b_net
  );
  bitbasher2 : entity xil_defaultlib.sysgen_bitbasher_086dfd1ec3 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in_x0 => fifo3_dout_net,
    a => bitbasher2_a_net,
    b => bitbasher2_b_net
  );
  bitbasher3 : entity xil_defaultlib.sysgen_bitbasher_086dfd1ec3 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in_x0 => fifo1_dout_net,
    a => bitbasher3_a_net,
    b => bitbasher3_b_net
  );
  bitbasher4 : entity xil_defaultlib.sysgen_bitbasher_086dfd1ec3 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in_x0 => fifo4_dout_net,
    a => bitbasher4_a_net,
    b => bitbasher4_b_net
  );
  bitbasher5 : entity xil_defaultlib.sysgen_bitbasher_086dfd1ec3 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in_x0 => fifo6_dout_net,
    a => bitbasher5_a_net,
    b => bitbasher5_b_net
  );
  bitbasher6 : entity xil_defaultlib.sysgen_bitbasher_086dfd1ec3 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in_x0 => fifo7_dout_net,
    a => bitbasher6_a_net,
    b => bitbasher6_b_net
  );
  bitbasher7 : entity xil_defaultlib.sysgen_bitbasher_086dfd1ec3 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in_x0 => fifo5_dout_net,
    a => bitbasher7_a_net,
    b => bitbasher7_b_net
  );
  bitbasher8 : entity xil_defaultlib.sysgen_bitbasher_086dfd1ec3 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in_x0 => fifo8_dout_net,
    a => bitbasher8_a_net,
    b => bitbasher8_b_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_71e89d757c 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net_x0
  );
  constant14 : entity xil_defaultlib.sysgen_constant_71e89d757c 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant14_op_net
  );
  constant15 : entity xil_defaultlib.sysgen_constant_a96178de4d 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant15_op_net
  );
  constant16 : entity xil_defaultlib.sysgen_constant_71e89d757c 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant16_op_net
  );
  constant2 : entity xil_defaultlib.sysgen_constant_71e89d757c 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant2_op_net_x0
  );
  constant3 : entity xil_defaultlib.sysgen_constant_71e89d757c 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant3_op_net_x0
  );
  constant4 : entity xil_defaultlib.sysgen_constant_71e89d757c 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant4_op_net_x0
  );
  constant5 : entity xil_defaultlib.sysgen_constant_71e89d757c 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant5_op_net_x0
  );
  constant6 : entity xil_defaultlib.sysgen_constant_71e89d757c 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant6_op_net_x0
  );
  delay1 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => gin_we_even_1_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay10 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => ts_6_net,
    clk => clk_net,
    ce => ce_net,
    q => delay10_q_net
  );
  delay11 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => ts_7_net,
    clk => clk_net,
    ce => ce_net,
    q => delay11_q_net_x0
  );
  delay12 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 8
  )
  port map (
    en => '1',
    rst => '0',
    d => ts_a_net,
    clk => clk_net,
    ce => ce_net,
    q => delay12_q_net
  );
  delay13 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 253,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => constant3_op_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay13_q_net
  );
  delay14 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => gin_tl_start_net,
    clk => clk_net,
    ce => ce_net,
    q => delay14_q_net
  );
  delay15 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay8_q_net_x3,
    clk => clk_net,
    ce => ce_net,
    q => delay15_q_net
  );
  delay16 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => ts_w_net,
    clk => clk_net,
    ce => ce_net,
    q => delay16_q_net
  );
  delay17 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 5,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay15_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay17_q_net
  );
  delay18 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 253,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => constant16_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay18_q_net
  );
  delay19 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d(0) => test_systolicfft_vhdl_black_box_vo_net,
    clk => clk_net,
    ce => ce_net,
    q => delay19_q_net
  );
  delay2 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => ts_0_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay26 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => gin_we_odd_2_net,
    clk => clk_net,
    ce => ce_net,
    q => delay26_q_net
  );
  delay28 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 253,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => constant14_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay28_q_net
  );
  delay29 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 253,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => constant2_op_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay29_q_net
  );
  delay3 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => ts_1_net,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  delay30 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 253,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => constant1_op_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay30_q_net
  );
  delay31 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => gin_we_even_3_net,
    clk => clk_net,
    ce => ce_net,
    q => delay31_q_net
  );
  delay35 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => gin_init_re_net,
    clk => clk_net,
    ce => ce_net,
    q => delay35_q_net
  );
  delay37 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 16
  )
  port map (
    en => '1',
    rst => '0',
    d => gin_dphi_net,
    clk => clk_net,
    ce => ce_net,
    q => delay37_q_net
  );
  delay38 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 8
  )
  port map (
    en => '1',
    rst => '0',
    d => gin_addr_net,
    clk => clk_net,
    ce => ce_net,
    q => delay38_q_net
  );
  delay4 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => ts_2_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net
  );
  delay43 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => gin_we_odd_4_net,
    clk => clk_net,
    ce => ce_net,
    q => delay43_q_net
  );
  delay44 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '0',
    d => gin_init_im_net,
    clk => clk_net,
    ce => ce_net,
    q => delay44_q_net
  );
  delay48 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => gin_we_odd_3_net,
    clk => clk_net,
    ce => ce_net,
    q => delay48_q_net
  );
  delay49 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => gin_we_even_4_net,
    clk => clk_net,
    ce => ce_net,
    q => delay49_q_net
  );
  delay5 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => ts_3_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  delay53 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 253,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => constant5_op_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay53_q_net
  );
  delay54 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 256,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => delay17_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay54_q_net
  );
  delay55 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 253,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => constant4_op_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay55_q_net
  );
  delay56 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 253,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => constant6_op_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay56_q_net
  );
  delay6 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => gin_we_odd_1_net,
    clk => clk_net,
    ce => ce_net,
    q => delay6_q_net
  );
  delay7 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => ts_4_net,
    clk => clk_net,
    ce => ce_net,
    q => delay7_q_net
  );
  delay8 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '0',
    d => gin_we_even_2_net,
    clk => clk_net,
    ce => ce_net,
    q => delay8_q_net
  );
  delay9 : entity xil_defaultlib.psb3_0_xldelay 
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 12
  )
  port map (
    en => '1',
    rst => '0',
    d => ts_5_net,
    clk => clk_net,
    ce => ce_net,
    q => delay9_q_net
  );
  expression : entity xil_defaultlib.sysgen_expr_dfc4963fbf 
  port map (
    clr => '0',
    a => register_q_net_x8,
    b => register_q_net_x9,
    clk => clk_net,
    ce => ce_net,
    dout => expression_dout_net
  );
  expression1 : entity xil_defaultlib.sysgen_expr_189d6fb430 
  port map (
    clr => '0',
    a1 => register_q_net_x2,
    a2 => register_q_net_x6,
    b1 => register_q_net_x1,
    b2 => register_q_net_x5,
    c1 => register_q_net_x0,
    c2 => register_q_net_x4,
    d1 => register_q_net,
    d2 => register_q_net_x3,
    clk => clk_net,
    ce => ce_net,
    dout => expression1_dout_net
  );
  fifo1 : entity xil_defaultlib.psb3_0_xlfifogen_u 
  generic map (
    core_name0 => "psb3_0_fifo_generator_i0",
    data_count_width => 10,
    data_width => 256,
    extra_registers => 1,
    has_ae => 0,
    has_af => 0,
    has_rst => false,
    ignore_din_for_gcd => false,
    percent_full_width => 1
  )
  port map (
    en => '1',
    rst => '0',
    din => concat1_y_net_x4,
    we => constant1_op_net_x0(0),
    re => delay30_q_net(0),
    clk => clk_net,
    ce => ce_net,
    we_ce => ce_net,
    re_ce => ce_net,
    dout => fifo1_dout_net,
    empty => fifo1_empty_net,
    full => fifo1_full_net
  );
  fifo2 : entity xil_defaultlib.psb3_0_xlfifogen_u 
  generic map (
    core_name0 => "psb3_0_fifo_generator_i0",
    data_count_width => 10,
    data_width => 256,
    extra_registers => 1,
    has_ae => 0,
    has_af => 0,
    has_rst => false,
    ignore_din_for_gcd => false,
    percent_full_width => 1
  )
  port map (
    en => '1',
    rst => '0',
    din => concat1_y_net_x6,
    we => constant14_op_net(0),
    re => delay28_q_net(0),
    clk => clk_net,
    ce => ce_net,
    we_ce => ce_net,
    re_ce => ce_net,
    dout => fifo2_dout_net,
    empty => fifo2_empty_net,
    full => fifo2_full_net
  );
  fifo3 : entity xil_defaultlib.psb3_0_xlfifogen_u 
  generic map (
    core_name0 => "psb3_0_fifo_generator_i0",
    data_count_width => 10,
    data_width => 256,
    extra_registers => 1,
    has_ae => 0,
    has_af => 0,
    has_rst => false,
    ignore_din_for_gcd => false,
    percent_full_width => 1
  )
  port map (
    en => '1',
    rst => '0',
    din => concat1_y_net_x5,
    we => constant16_op_net(0),
    re => delay18_q_net(0),
    clk => clk_net,
    ce => ce_net,
    we_ce => ce_net,
    re_ce => ce_net,
    dout => fifo3_dout_net,
    empty => fifo3_empty_net,
    full => fifo3_full_net
  );
  fifo4 : entity xil_defaultlib.psb3_0_xlfifogen_u 
  generic map (
    core_name0 => "psb3_0_fifo_generator_i0",
    data_count_width => 10,
    data_width => 256,
    extra_registers => 1,
    has_ae => 0,
    has_af => 0,
    has_rst => false,
    ignore_din_for_gcd => false,
    percent_full_width => 1
  )
  port map (
    en => '1',
    rst => '0',
    din => concat1_y_net_x3,
    we => constant2_op_net_x0(0),
    re => delay29_q_net(0),
    clk => clk_net,
    ce => ce_net,
    we_ce => ce_net,
    re_ce => ce_net,
    dout => fifo4_dout_net,
    empty => fifo4_empty_net,
    full => fifo4_full_net
  );
  fifo5 : entity xil_defaultlib.psb3_0_xlfifogen_u 
  generic map (
    core_name0 => "psb3_0_fifo_generator_i0",
    data_count_width => 10,
    data_width => 256,
    extra_registers => 1,
    has_ae => 0,
    has_af => 0,
    has_rst => false,
    ignore_din_for_gcd => false,
    percent_full_width => 1
  )
  port map (
    en => '1',
    rst => '0',
    din => concat1_y_net_x0,
    we => constant3_op_net_x0(0),
    re => delay13_q_net(0),
    clk => clk_net,
    ce => ce_net,
    we_ce => ce_net,
    re_ce => ce_net,
    dout => fifo5_dout_net,
    empty => fifo5_empty_net,
    full => fifo5_full_net
  );
  fifo6 : entity xil_defaultlib.psb3_0_xlfifogen_u 
  generic map (
    core_name0 => "psb3_0_fifo_generator_i0",
    data_count_width => 10,
    data_width => 256,
    extra_registers => 1,
    has_ae => 0,
    has_af => 0,
    has_rst => false,
    ignore_din_for_gcd => false,
    percent_full_width => 1
  )
  port map (
    en => '1',
    rst => '0',
    din => concat1_y_net_x2,
    we => constant4_op_net_x0(0),
    re => delay55_q_net(0),
    clk => clk_net,
    ce => ce_net,
    we_ce => ce_net,
    re_ce => ce_net,
    dout => fifo6_dout_net,
    empty => fifo6_empty_net,
    full => fifo6_full_net
  );
  fifo7 : entity xil_defaultlib.psb3_0_xlfifogen_u 
  generic map (
    core_name0 => "psb3_0_fifo_generator_i0",
    data_count_width => 10,
    data_width => 256,
    extra_registers => 1,
    has_ae => 0,
    has_af => 0,
    has_rst => false,
    ignore_din_for_gcd => false,
    percent_full_width => 1
  )
  port map (
    en => '1',
    rst => '0',
    din => concat1_y_net_x1,
    we => constant5_op_net_x0(0),
    re => delay53_q_net(0),
    clk => clk_net,
    ce => ce_net,
    we_ce => ce_net,
    re_ce => ce_net,
    dout => fifo7_dout_net,
    empty => fifo7_empty_net,
    full => fifo7_full_net
  );
  fifo8 : entity xil_defaultlib.psb3_0_xlfifogen_u 
  generic map (
    core_name0 => "psb3_0_fifo_generator_i0",
    data_count_width => 10,
    data_width => 256,
    extra_registers => 1,
    has_ae => 0,
    has_af => 0,
    has_rst => false,
    ignore_din_for_gcd => false,
    percent_full_width => 1
  )
  port map (
    en => '1',
    rst => '0',
    din => concat1_y_net,
    we => constant6_op_net_x0(0),
    re => delay56_q_net(0),
    clk => clk_net,
    ce => ce_net,
    we_ce => ce_net,
    re_ce => ce_net,
    dout => fifo8_dout_net,
    empty => fifo8_empty_net,
    full => fifo8_full_net
  );
  ram_dphi_addr : entity xil_defaultlib.psb3_0_xlcounter_free 
  generic map (
    core_name0 => "psb3_0_c_counter_binary_v12_0_i0",
    op_arith => xlUnsigned,
    op_width => 8
  )
  port map (
    clr => '0',
    rst => gin_tl_reset_net,
    en => gin_tl_start_net,
    clk => clk_net,
    ce => ce_net,
    op => ram_dphi_addr_op_net
  );
  reinterpret : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => bitbasher1_b_net,
    output_port => reinterpret_output_port_net
  );
  reinterpret1 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => bitbasher3_b_net,
    output_port => reinterpret1_output_port_net_x14
  );
  reinterpret2 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => bitbasher4_b_net,
    output_port => reinterpret2_output_port_net_x14
  );
  reinterpret3 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => bitbasher2_b_net,
    output_port => reinterpret3_output_port_net_x14
  );
  reinterpret4 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => bitbasher5_b_net,
    output_port => reinterpret4_output_port_net_x14
  );
  reinterpret5 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => bitbasher7_b_net,
    output_port => reinterpret5_output_port_net_x14
  );
  reinterpret6 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => bitbasher8_b_net,
    output_port => reinterpret6_output_port_net_x14
  );
  reinterpret7 : entity xil_defaultlib.sysgen_reinterpret_5672cd6a95 
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => bitbasher6_b_net,
    output_port => reinterpret7_output_port_net_x14
  );
end structural;
-- Generated from Simulink block 
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0_default_clock_driver is
  port (
    psb3_0_sysclk : in std_logic;
    psb3_0_sysce : in std_logic;
    psb3_0_sysclr : in std_logic;
    psb3_0_clk1 : out std_logic;
    psb3_0_ce1 : out std_logic
  );
end psb3_0_default_clock_driver;
architecture structural of psb3_0_default_clock_driver is 
begin
  clockdriver : entity xil_defaultlib.xlclockdriver 
  generic map (
    period => 1,
    log_2_period => 1
  )
  port map (
    sysclk => psb3_0_sysclk,
    sysce => psb3_0_sysce,
    sysclr => psb3_0_sysclr,
    clk => psb3_0_clk1,
    ce => psb3_0_ce1
  );
end structural;
-- Generated from Simulink block 
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity psb3_0 is
  port (
    gin_tl_reset : in std_logic_vector( 1-1 downto 0 );
    gin_tl_start : in std_logic_vector( 1-1 downto 0 );
    gin_addr : in std_logic_vector( 8-1 downto 0 );
    gin_dphi : in std_logic_vector( 16-1 downto 0 );
    gin_init_im : in std_logic_vector( 18-1 downto 0 );
    gin_init_re : in std_logic_vector( 18-1 downto 0 );
    gin_we_even_1 : in std_logic_vector( 1-1 downto 0 );
    gin_we_even_2 : in std_logic_vector( 1-1 downto 0 );
    gin_we_even_3 : in std_logic_vector( 1-1 downto 0 );
    gin_we_even_4 : in std_logic_vector( 1-1 downto 0 );
    gin_we_odd_1 : in std_logic_vector( 1-1 downto 0 );
    gin_we_odd_2 : in std_logic_vector( 1-1 downto 0 );
    gin_we_odd_3 : in std_logic_vector( 1-1 downto 0 );
    gin_we_odd_4 : in std_logic_vector( 1-1 downto 0 );
    ts_0 : in std_logic_vector( 12-1 downto 0 );
    ts_1 : in std_logic_vector( 12-1 downto 0 );
    ts_2 : in std_logic_vector( 12-1 downto 0 );
    ts_3 : in std_logic_vector( 12-1 downto 0 );
    ts_4 : in std_logic_vector( 12-1 downto 0 );
    ts_5 : in std_logic_vector( 12-1 downto 0 );
    ts_6 : in std_logic_vector( 12-1 downto 0 );
    ts_7 : in std_logic_vector( 12-1 downto 0 );
    ts_a : in std_logic_vector( 8-1 downto 0 );
    ts_w : in std_logic_vector( 1-1 downto 0 );
    clk : in std_logic;
    gout_cordic_delay_even_1 : out std_logic_vector( 12-1 downto 0 );
    gout_psb_tvalid : out std_logic_vector( 1-1 downto 0 );
    gout_delay_ifft : out std_logic_vector( 12-1 downto 0 );
    gout_ov_ifft : out std_logic_vector( 1-1 downto 0 );
    gout_ov_add : out std_logic_vector( 1-1 downto 0 );
    gout_psb_im_0 : out std_logic_vector( 16-1 downto 0 );
    gout_psb_im_1 : out std_logic_vector( 16-1 downto 0 );
    gout_psb_im_2 : out std_logic_vector( 16-1 downto 0 );
    gout_psb_im_3 : out std_logic_vector( 16-1 downto 0 );
    gout_psb_re_0 : out std_logic_vector( 16-1 downto 0 );
    gout_psb_re_1 : out std_logic_vector( 16-1 downto 0 );
    gout_psb_re_2 : out std_logic_vector( 16-1 downto 0 );
    gout_psb_re_3 : out std_logic_vector( 16-1 downto 0 )
  );
end psb3_0;
architecture structural of psb3_0 is 
  attribute core_generation_info : string;
  attribute core_generation_info of structural : architecture is "psb3_0,sysgen_core_2021_1,{,compilation=IP Catalog,block_icon_display=Default,family=zynquplusRFSOC,part=xczu28dr,speed=-2-e,package=ffvg1517,synthesis_language=vhdl,hdl_library=xil_defaultlib,synthesis_strategy=Vivado Synthesis Defaults,implementation_strategy=Vivado Implementation Defaults,testbench=0,interface_doc=1,ce_clr=0,clock_period=10,system_simulink_period=1,waveform_viewer=0,axilite_interface=0,ip_catalog_plugin=0,hwcosim_burst_mode=0,simulation_time=3000,abs=32,accum=1,addsub=152,bitbasher=48,blackbox2=1,concat=42,constant=163,convert=17,cordic_v6_0=8,counter=48,delay=460,dpram=44,expr=12,fifo=32,inv=9,logical=17,mult=128,mux=129,register=45,reinterpret=544,relational=34,slice=880,spram=32,}";
  signal clk_1_net : std_logic;
  signal ce_1_net : std_logic;
begin
  psb3_0_default_clock_driver : entity xil_defaultlib.psb3_0_default_clock_driver 
  port map (
    psb3_0_sysclk => clk,
    psb3_0_sysce => '1',
    psb3_0_sysclr => '0',
    psb3_0_clk1 => clk_1_net,
    psb3_0_ce1 => ce_1_net
  );
  psb3_0_struct : entity xil_defaultlib.psb3_0_struct 
  port map (
    gin_tl_reset => gin_tl_reset,
    gin_tl_start => gin_tl_start,
    gin_addr => gin_addr,
    gin_dphi => gin_dphi,
    gin_init_im => gin_init_im,
    gin_init_re => gin_init_re,
    gin_we_even_1 => gin_we_even_1,
    gin_we_even_2 => gin_we_even_2,
    gin_we_even_3 => gin_we_even_3,
    gin_we_even_4 => gin_we_even_4,
    gin_we_odd_1 => gin_we_odd_1,
    gin_we_odd_2 => gin_we_odd_2,
    gin_we_odd_3 => gin_we_odd_3,
    gin_we_odd_4 => gin_we_odd_4,
    ts_0 => ts_0,
    ts_1 => ts_1,
    ts_2 => ts_2,
    ts_3 => ts_3,
    ts_4 => ts_4,
    ts_5 => ts_5,
    ts_6 => ts_6,
    ts_7 => ts_7,
    ts_a => ts_a,
    ts_w => ts_w,
    clk_1 => clk_1_net,
    ce_1 => ce_1_net,
    gout_cordic_delay_even_1 => gout_cordic_delay_even_1,
    gout_psb_tvalid => gout_psb_tvalid,
    gout_delay_ifft => gout_delay_ifft,
    gout_ov_ifft => gout_ov_ifft,
    gout_ov_add => gout_ov_add,
    gout_psb_im_0 => gout_psb_im_0,
    gout_psb_im_1 => gout_psb_im_1,
    gout_psb_im_2 => gout_psb_im_2,
    gout_psb_im_3 => gout_psb_im_3,
    gout_psb_re_0 => gout_psb_re_0,
    gout_psb_re_1 => gout_psb_re_1,
    gout_psb_re_2 => gout_psb_re_2,
    gout_psb_re_3 => gout_psb_re_3
  );
end structural;
